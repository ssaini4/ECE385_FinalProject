module font_poke ( input [8:0] addr, output [23:0] data);
					 
parameter DATA_WIDTH = 24;

parameter [0:899][DATA_WIDTH-1:0] poke = {
24'hffffff, 24'hffffff, 24'hffffff, 24'hffffff, 24'hffffff, 24'hffffff, 24'hffffff, 24'hffffff, 24'hffffff, 24'hffffff, 24'hffffff, 24'hffffff, 24'hffffff, 24'hffffff, 24'hffffff, 24'hffffff, 24'hffffff, 24'hffffff, 24'hffffff, 24'h000, 24'h000, 24'hffffff, 24'hffffff, 24'hffffff, 24'hffffff, 24'hffffff, 24'hffffff, 24'hffffff, 24'hffffff, 24'hffffff, 24'hffffff, 24'h000, 24'h000, 24'h000, 24'h000, 24'hffffff, 24'hffffff, 24'hffffff, 24'hffffff, 24'hffffff, 24'hffffff, 24'hffffff, 24'hffffff, 24'hffffff, 24'hffffff, 24'hffffff, 24'hffffff, 24'hffffff, 24'h111, 24'h000, 24'h000, 24'hffffff, 24'hffffff, 24'hffffff, 24'hffffff, 24'hffffff, 24'hffffff, 24'hffffff, 24'hffffff, 24'hffffff, 24'hffffff, 24'hffffff, 24'h000, 24'h000, 24'h000, 24'h000, 24'h000, 24'hffffff, 24'hffffff, 24'hffffff, 24'hffffff, 24'hffffff, 24'hffffff, 24'hffffff, 24'hffffff, 24'hffffff, 24'hffffff, 24'h444, 24'h000, 24'h000, 24'h000, 24'hffffff, 24'hffffff, 24'hffffff, 24'hffffff, 24'hffffff, 24'hffffff, 24'hffffff, 24'hffffff, 24'hffffff, 24'hffffff, 24'hffffff, 24'hffffff, 24'h000, 24'h000, 24'hf0c516, 24'hf0c516, 24'h161b15, 24'h000, 24'hffffff, 24'hffffff, 24'hffffff, 24'hffffff, 24'hffffff, 24'hffffff, 24'hffffff, 24'hffffff, 24'h000, 24'hf7c21e, 24'h024, 24'h000, 24'hffffff, 24'hffffff, 24'hffffff, 24'hffffff, 24'hffffff, 24'hffffff, 24'hffffff, 24'hffffff, 24'hffffff, 24'hffffff, 24'hffffff, 24'hffffff, 24'hffffff, 24'h000, 24'hd3a12, 24'hf6c31a, 24'he9c332, 24'hc50, 24'h000, 24'h000, 24'hffffff, 24'hffffff, 24'hffffff, 24'hffffff, 24'hffffff, 24'h000, 24'hf7c121, 24'hf7c510, 24'h602, 24'h000, 24'hffffff, 24'hffffff, 24'hffffff, 24'hffffff, 24'hffffff, 24'hffffff, 24'hffffff, 24'hffffff, 24'hffffff, 24'hffffff, 24'hffffff, 24'hffffff, 24'hffffff, 24'hffffff, 24'h02b, 24'hd39d0, 24'hf6c31c, 24'hf3c227, 24'hefc9e, 24'he1c74c, 24'h000, 24'h000, 24'h000, 24'h000, 24'hffffff, 24'h000, 24'hf6c31c, 24'hf7c41b, 24'h602, 24'hffffff, 24'hffffff, 24'hffffff, 24'hffffff, 24'hffffff, 24'hffffff, 24'hffffff, 24'hffffff, 24'hffffff, 24'hffffff, 24'hffffff, 24'hffffff, 24'hffffff, 24'hffffff, 24'hffffff, 24'h000, 24'hd2a00, 24'hf6c318, 24'hf6c417, 24'hf6c31c, 24'he9c316, 24'he2c454, 24'he2c454, 24'he2c454, 24'he2c454, 24'h000, 24'h000, 24'hf6c31c, 24'hd09e0, 24'h600, 24'hffffff, 24'hffffff, 24'hffffff, 24'hffffff, 24'hffffff, 24'hffffff, 24'hffffff, 24'hffffff, 24'hffffff, 24'hffffff, 24'hffffff, 24'hffffff, 24'hffffff, 24'hffffff, 24'hffffff, 24'hffffff, 24'h000, 24'h000, 24'he3c360, 24'hf6c31c, 24'hf6c31c, 24'hf6c31c, 24'hf6c31c, 24'hf6c31c, 24'hf6c31c, 24'h027, 24'h027, 24'hf6c31c, 24'hd09e0, 24'h600, 24'hffffff, 24'hffffff, 24'hffffff, 24'hffffff, 24'hffffff, 24'hffffff, 24'hffffff, 24'hffffff, 24'hffffff, 24'hffffff, 24'hffffff, 24'hffffff, 24'hffffff, 24'hffffff, 24'hffffff, 24'hffffff, 24'hffffff, 24'h000, 24'hdcbf6f, 24'heac435, 24'he9c732, 24'hf6c31c, 24'hf6c31c, 24'hf6c31c, 24'hf6c31c, 24'hf6c31c, 24'hf6c31c, 24'hf6c31c, 24'hc69e22, 24'h030, 24'hffffff, 24'hffffff, 24'hffffff, 24'hffffff, 24'hffffff, 24'hffffff, 24'hffffff, 24'hffffff, 24'hffffff, 24'hffffff, 24'hffffff, 24'hffffff, 24'hffffff, 24'hffffff, 24'hffffff, 24'hffffff, 24'hffffff, 24'h0e0, 24'h700, 24'h000, 24'hfff9ff, 24'hf6c31c, 24'hf6c31c, 24'hf6c31c, 24'hf6c31c, 24'hf6c31c, 24'hf6c31c, 24'hf6c31c, 24'h300, 24'hffffff, 24'hffffff, 24'hffffff, 24'hffffff, 24'hffffff, 24'hffffff, 24'hffffff, 24'hffffff, 24'hffffff, 24'hffffff, 24'hffffff, 24'hffffff, 24'hffffff, 24'hffffff, 24'hffffff, 24'hffffff, 24'hffffff, 24'h1b00, 24'he30b, 24'h4500, 24'h012, 24'h00b, 24'hf6c31c, 24'hf6c31c, 24'hf6c31c, 24'hf6c31c, 24'hf3c26, 24'hfac9d, 24'hf6c31c, 24'h300, 24'hffffff, 24'hffffff, 24'hffffff, 24'hffffff, 24'hffffff, 24'hffffff, 24'hffffff, 24'hffffff, 24'hffffff, 24'hffffff, 24'hffffff, 24'hffffff, 24'hffffff, 24'hffffff, 24'hffffff, 24'hffffff, 24'h000, 24'hd137, 24'hdc00, 24'hffa53d, 24'hf6c31c, 24'hf6c31c, 24'hf6c31c, 24'hf6c31c, 24'hf6c31c, 24'hf6c31c, 24'hffffff, 24'h000, 24'hf6c31c, 24'h300, 24'hffffff, 24'hffffff, 24'hffffff, 24'hffffff, 24'hffffff, 24'hffffff, 24'hffffff, 24'hffffff, 24'hffffff, 24'hffffff, 24'hffffff, 24'hffffff, 24'hffffff, 24'hffffff, 24'hffffff, 24'hffffff, 24'h000, 24'hbee0, 24'hd920, 24'hffa53d, 24'hf6c31c, 24'hf6c31c, 24'hf6c31c, 24'hf6c31c, 24'hf6c31c, 24'hf6c31c, 24'h304, 24'he00, 24'hf4c41a, 24'h020, 24'hffffff, 24'hffffff, 24'hffffff, 24'hffffff, 24'hffffff, 24'hffffff, 24'hffffff, 24'hffffff, 24'hffffff, 24'hffffff, 24'hffffff, 24'hffffff, 24'hffffff, 24'hffffff, 24'hffffff, 24'hffffff, 24'hffffff, 24'h000, 24'hf000, 24'hffa53d, 24'hf6c31c, 24'hf6c31c, 24'hf6c31c, 24'hf6c31c, 24'hf6c31c, 24'hf6c31c, 24'hf6c31c, 24'hdc00, 24'h000, 24'h000, 24'h000, 24'h000, 24'hffffff, 24'hffffff, 24'hffffff, 24'hffffff, 24'hffffff, 24'hffffff, 24'hffffff, 24'hffffff, 24'hffffff, 24'hffffff, 24'hffffff, 24'hffffff, 24'hffffff, 24'hffffff, 24'h000, 24'h000, 24'h000, 24'h000, 24'h040, 24'hf6c31c, 24'hf6c31c, 24'hf6c31c, 24'hf6c31c, 24'hf6c31c, 24'hdc00, 24'hdc00, 24'h000, 24'hf8c21a, 24'hf6c31c, 24'hf6c31c, 24'h607, 24'h222, 24'hffffff, 24'hffffff, 24'hffffff, 24'hffffff, 24'hffffff, 24'hffffff, 24'hffffff, 24'hffffff, 24'hffffff, 24'hffffff, 24'hffffff, 24'h000, 24'hf6c31c, 24'hf6c31c, 24'hf6c31c, 24'hf6c31c, 24'hfabf23, 24'h002, 24'hf6c31c, 24'hf6c31c, 24'hf6c31c, 24'hf6c31c, 24'hdc00, 24'h000, 24'hf6c31c, 24'hf6c31c, 24'hf6c31c, 24'h304, 24'h000, 24'h000, 24'h000, 24'h000, 24'h000, 24'h000, 24'hffffff, 24'hffffff, 24'hffffff, 24'hffffff, 24'hffffff, 24'hffffff, 24'h000, 24'hf6c31c, 24'hf6c31c, 24'hf6c31c, 24'hf6c31c, 24'hf6c31c, 24'hf6c31c, 24'hfac118, 24'h300, 24'hd09e1, 24'hf6c31c, 24'hf6c31c, 24'h000, 24'hf6c31c, 24'hf6c31c, 24'hcda00, 24'h307, 24'hfabf23, 24'hf6c31c, 24'hf6c31c, 24'hf6c31c, 24'hf6c31c, 24'hf6c31c, 24'hf6c31c, 24'h000, 24'h000, 24'h000, 24'hffffff, 24'hffffff, 24'hffffff, 24'hffffff, 24'h000, 24'hd09e1, 24'hd09e1, 24'hd09e1, 24'hd09e1, 24'hd09e1, 24'hd09e0, 24'h600, 24'hf6c31c, 24'hf6c31c, 24'hf6c31c, 24'hf6c31c, 24'hf6c31c, 24'hd09e1, 24'h104, 24'hefc61c, 24'hd09d3, 24'hf8c724, 24'hf6c31c, 24'hf6c31c, 24'hf6c31c, 24'hf6c31c, 24'hf6c31c, 24'hf6c31c, 24'hf6c31c, 24'hf6c31c, 24'hffffff, 24'hffffff, 24'hffffff, 24'hffffff, 24'hffffff, 24'h000, 24'h000, 24'h000, 24'h000, 24'h000, 24'h002, 24'hf6c31c, 24'hf6c31c, 24'hf6c31c, 24'hf6c31c, 24'hf6c31c, 24'hd09e1, 24'h000, 24'h000, 24'hefc61c, 24'hd09d3, 24'hd09e1, 24'hf6c31c, 24'hf6c31c, 24'hf6c31c, 24'hf6c31c, 24'hf6c31c, 24'hf6c31c, 24'hf6c31c, 24'h000, 24'hffffff, 24'hffffff, 24'hffffff, 24'hffffff, 24'hffffff, 24'h000, 24'hf5bb1c, 24'hf6c31c, 24'hf6c31c, 24'hf6c31c, 24'hf6c31c, 24'hf6c31c, 24'hf6c31c, 24'hf6c31c, 24'hf6c31c, 24'hf6c31c, 24'h000, 24'hffffff, 24'h000, 24'hefc61c, 24'hd09d3, 24'hd09e1, 24'hd09e1, 24'hd09e1, 24'hcf9d0, 24'hf6c31c, 24'hf6c31c, 24'hf6c31c, 24'h000, 24'hffffff, 24'hffffff, 24'hffffff, 24'hffffff, 24'hffffff, 24'hffffff, 24'h000, 24'hf5bb1c, 24'hf6c31c, 24'hf6c31c, 24'hf6c31c, 24'hf6c31c, 24'hf6c31c, 24'hf6c31c, 24'hf6c31c, 24'hf6c31c, 24'hf6c31c, 24'h000, 24'h000, 24'h000, 24'hefc61c, 24'hd09d3, 24'h1500, 24'h000, 24'h000, 24'hf00, 24'hd09e1, 24'hf6c31c, 24'h000, 24'hffffff, 24'hffffff, 24'hffffff, 24'hffffff, 24'hffffff, 24'hffffff, 24'h000, 24'hf6c31c, 24'hf6c31c, 24'hf6c31c, 24'hf6c31c, 24'hf6c31c, 24'hf6c31c, 24'hf6c31c, 24'hf6c31c, 24'hf6c31c, 24'hf6c31c, 24'hf6c31c, 24'h000, 24'hd09e1, 24'hd09e1, 24'hd09e1, 24'h001b, 24'hffffff, 24'hffffff, 24'hffffff, 24'hfcfcfc, 24'h000, 24'h000, 24'hffffff, 24'hffffff, 24'hffffff, 24'hffffff, 24'hffffff, 24'hffffff, 24'hffffff, 24'h000, 24'hf6c31c, 24'hf6c31c, 24'hf6c31c, 24'hf6c31c, 24'hf6c31c, 24'hf6c31c, 24'hf6c31c, 24'hf6c31c, 24'hf6c31c, 24'hf6c31c, 24'hf6c31c, 24'h000, 24'h72281, 24'h100, 24'h000, 24'hffffff, 24'hffffff, 24'hffffff, 24'hffffff, 24'hffffff, 24'hffffff, 24'hffffff, 24'hffffff, 24'hffffff, 24'hffffff, 24'hffffff, 24'hffffff, 24'hffffff, 24'h000, 24'hf6c31c, 24'hf6c31c, 24'hf6c31c, 24'hf6c31c, 24'hf6c31c, 24'hf6c31c, 24'hf6c31c, 24'hf6c31c, 24'hf6c31c, 24'hf6c31c, 24'hf6c31c, 24'hf6c31c, 24'h72281, 24'h72281, 24'h100, 24'hffffff, 24'hffffff, 24'hffffff, 24'hffffff, 24'hffffff, 24'hffffff, 24'hffffff, 24'hffffff, 24'hffffff, 24'hffffff, 24'hffffff, 24'hffffff, 24'hffffff, 24'hffffff, 24'h000, 24'hd09e1, 24'hd09e1, 24'hf8c51e, 24'hf6c31c, 24'hf6c31c, 24'hf6c31c, 24'hf6c31c, 24'hf6c31c, 24'hf6c31c, 24'hf6c31c, 24'hf6c31c, 24'hf6c31c, 24'hf6c31c, 24'h000, 24'hffffff, 24'hffffff, 24'hffffff, 24'hffffff, 24'hffffff, 24'hffffff, 24'hffffff, 24'hffffff, 24'hffffff, 24'hffffff, 24'hffffff, 24'hffffff, 24'hffffff, 24'hffffff, 24'hffffff, 24'hffffff, 24'h000, 24'hd09e1, 24'hd09e1, 24'hd09e1, 24'hd09e1, 24'hd09e1, 24'hd09e1, 24'hd09e1, 24'hd09e1, 24'hd09e1, 24'hd09e1, 24'hf6c31c, 24'h000, 24'hffffff, 24'hffffff, 24'hffffff, 24'hffffff, 24'hffffff, 24'hffffff, 24'hffffff, 24'hffffff, 24'hffffff, 24'hffffff, 24'hffffff, 24'hffffff, 24'hffffff, 24'hffffff, 24'hffffff, 24'hffffff, 24'h000, 24'hfebe1e, 24'hd09e1, 24'hd09e1, 24'hf0b, 24'h090, 24'h090, 24'h090, 24'h090, 24'h090, 24'h090, 24'hd09e1, 24'hd09e0, 24'hfabd2f, 24'h000, 24'hffffff, 24'hffffff, 24'hffffff, 24'hffffff, 24'hffffff, 24'hffffff, 24'hffffff, 24'hffffff, 24'hffffff, 24'hffffff, 24'hffffff, 24'hffffff, 24'hffffff, 24'hffffff, 24'hffffff, 24'hffffff, 24'h012, 24'h100, 24'h100, 24'hfeffff, 24'hffffff, 24'hffffff, 24'hffffff, 24'hffffff, 24'hffffff, 24'hffffff, 24'h100, 24'h100, 24'hf6c31c, 24'hf3c41e, 24'h304, 24'hffffff, 24'hffffff, 24'hffffff, 24'hffffff, 24'hffffff, 24'hffffff, 24'hffffff, 24'hffffff, 24'hffffff, 24'hffffff, 24'hffffff, 24'hffffff, 24'hffffff, 24'hffffff, 24'hffffff, 24'hffffff, 24'hffffff, 24'hffffff, 24'hffffff, 24'hffffff, 24'hffffff, 24'hffffff, 24'hffffff, 24'hffffff, 24'hffffff, 24'hffffff, 24'hffffff, 24'h300, 24'h300, 24'hfffeff, 24'hffffff, 24'hffffff, 24'hffffff, 24'hffffff, 24'hffffff, 24'hffffff, 24'hffffff, 24'hffffff, 24'hffffff, 24'hffffff, 24'hffffff, 24'hfffdf3, 24'hfffdf3, 24'hfffdf3, 24'hfffdf3, 24'hfffdf3, 24'hfffdf3, 24'hfffdf3, 24'hfffdf3, 24'hfffdf3, 24'hfffdf3, 24'hfffdf3, 24'hfffdf3, 24'hfffdf3, 24'hfffdf3, 24'hfffdf3, 24'hfffdf3, 24'hfffdf3, 24'hfffdf3, 24'hfffdf3, 24'hfffdf3, 24'hfffdf3, 24'hfffdf3, 24'hfffdf3, 24'hfffdf3, 24'hfffdf3, 24'hfffdf3, 24'hfffdf3, 24'hfffdf3, 24'hfffdf3, 24'hfffdf3
};
assign data = poke[addr];

endmodule
