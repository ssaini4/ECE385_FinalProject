module font_start ( input [19:0] addr, output [7:0] data);
					 
parameter DATA_WIDTH = 8;
parameter [0:510*210-1][DATA_WIDTH-1:0] screen = {8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h1a,8'h1a,8'h1a,8'h1a,8'h1a,8'h1a,8'h1a,8'h1a,8'h1a,8'h1a,8'h1a,8'h1a,8'h1a,8'h1a,8'h1a,8'h1a,8'h2b,8'h1a,8'h1a,8'h1a,8'h1a,8'h1a,8'h2b,8'h1a,8'h1a,8'h2b,8'h1a,8'h1a,8'h1a,8'h1a,8'h1a,8'h1a,8'h1a,8'h1a,8'h1a,8'h1a,8'h1a,8'h1a,8'h1a,8'h1a,8'h1a,8'h1a,8'h1a,8'h1a,8'h1a,8'h1a,8'h1a,8'h1a,8'h1a,8'h2b,8'h1a,8'h2b,8'h1a,8'h1a,8'h1a,8'h1a,8'h2b,8'h1a,8'h1a,8'h1a,8'h1a,8'h1a,8'h2b,8'h1a,8'h1a,8'h1a,8'h1a,8'h1a,8'h1a,8'h1a,8'h1a,8'h1a,8'h1a,8'h1a,8'h2b,8'h2b,8'h1a,8'h1a,8'h2b,8'h2b,8'h2b,8'h1a,8'h1a,8'h1a,8'h1a,8'h1a,8'h1a,8'h2b,8'h1a,8'h1a,8'h1a,8'h1a,8'h1a,8'h1a,8'h1a,8'h1a,8'h1a,8'h1a,8'h1a,8'h2b,8'h1a,8'h1a,8'h2b,8'h1a,8'h1a,8'h1a,8'h2b,8'h1a,8'h1a,8'h1a,8'h1a,8'h1a,8'h2b,8'h1a,8'h1a,8'h2b,8'h1a,8'h1a,8'h1a,8'h1a,8'h1a,8'h1a,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h1a,8'h1a,8'h1a,8'h1a,8'h1a,8'h1a,8'h2b,8'h2b,8'h1a,8'h1a,8'h1a,8'h1a,8'h1a,8'h1a,8'h1a,8'h1a,8'h2b,8'h2b,8'h1a,8'h1a,8'h1a,8'h1a,8'h1a,8'h1a,8'h1a,8'h2b,8'h2b,8'h1a,8'h1a,8'h1a,8'h1a,8'h1a,8'h1a,8'h1a,8'h1a,8'h1a,8'h1a,8'h1a,8'h1a,8'h1a,8'h2b,8'h1a,8'h1a,8'h1a,8'h1a,8'h1a,8'h1a,8'h1a,8'h2b,8'h2b,8'h1a,8'h1a,8'h1a,8'h1a,8'h1a,8'h1a,8'h1a,8'h2b,8'h1a,8'h1a,8'h1a,8'h1a,8'h1a,8'h2b,8'h2b,8'h2b,8'h1a,8'h1a,8'h1a,8'h1a,8'h1a,8'h1a,8'h1a,8'h1a,8'h2b,8'h2b,8'h1a,8'h1a,8'h1a,8'h1a,8'h1a,8'h1a,8'h1a,8'h1a,8'h2b,8'h1a,8'h1a,8'h1a,8'h1a,8'h1a,8'h1a,8'h1a,8'h1a,8'h1a,8'h1a,8'h1a,8'h1a,8'h2b,8'h2b,8'h2b,8'h1a,8'h1a,8'h1a,8'h1a,8'h1a,8'h1a,8'h1a,8'h1a,8'h1a,8'h1a,8'h1a,8'h1a,8'h1a,8'h2b,8'h2b,8'h2b,8'h1a,8'h1a,8'h1a,8'h1a,8'h1a,8'h1a,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h1a,8'h1a,8'h1a,8'h1a,8'h1a,8'h1a,8'h1a,8'h1a,8'h1a,8'h1a,8'h1a,8'h1a,8'h1a,8'h1a,8'h1a,8'h1a,8'h1a,8'h2b,8'h1a,8'h1a,8'h1a,8'h21,8'h6,8'h9,8'h2b,8'h1a,8'h1a,8'h1a,8'h1a,8'h1a,8'h2b,8'h1a,8'h1a,8'h2b,8'h1a,8'h1a,8'h1a,8'h1a,8'h2b,8'h2b,8'h1a,8'h1a,8'h1a,8'h1a,8'h1a,8'h1a,8'h2b,8'h1a,8'h2b,8'h1a,8'h1a,8'h2b,8'h1a,8'h1a,8'h1a,8'h1a,8'h2b,8'h2b,8'h1a,8'h1a,8'h2b,8'h2b,8'h1a,8'h1a,8'h1a,8'h1a,8'h1a,8'h1a,8'h1a,8'h1a,8'h2b,8'h1a,8'h1a,8'h1a,8'h1a,8'h1a,8'h1a,8'h1a,8'h1a,8'h1a,8'h1a,8'h2b,8'h1a,8'h1a,8'h1a,8'h2b,8'h1a,8'h1a,8'h1a,8'h1a,8'h1a,8'h2b,8'h2b,8'h2b,8'h1a,8'h1a,8'h1a,8'h2b,8'h1a,8'h1a,8'h1a,8'h2b,8'h2b,8'h1a,8'h2b,8'h1a,8'h1a,8'h1a,8'h2b,8'h2b,8'h2b,8'h2b,8'h1a,8'h2b,8'h2b,8'h1a,8'h1a,8'h2b,8'h1a,8'h1a,8'h1a,8'h1a,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h1a,8'h21,8'h6,8'h6,8'h6,8'h6,8'h6,8'h6,8'h1b,8'h1a,8'h1a,8'h1a,8'h1a,8'h1a,8'h1a,8'h1a,8'h1a,8'h2b,8'h1a,8'h1a,8'h1a,8'h21,8'h6,8'h22,8'h1a,8'h1a,8'h2b,8'h1a,8'h1a,8'h1a,8'h1a,8'h1a,8'h1a,8'h2b,8'h1a,8'h2b,8'h2b,8'h1a,8'h1a,8'h2b,8'h1a,8'h1a,8'h1a,8'h1a,8'h1a,8'h1a,8'h1a,8'h1a,8'h1a,8'h1a,8'h1a,8'h2b,8'h1a,8'h1a,8'h1a,8'h1a,8'h1a,8'h1a,8'h1a,8'h1a,8'h2b,8'h1a,8'h2b,8'h2b,8'h1a,8'h1a,8'h1a,8'h2b,8'h1a,8'h1a,8'h2b,8'h1a,8'h1a,8'h1a,8'h1a,8'h1a,8'h1a,8'h1a,8'h1a,8'h1a,8'h1a,8'h6,8'h6,8'h6,8'h6,8'h6,8'h2a,8'h1a,8'h1a,8'h1a,8'h1a,8'h1a,8'h22,8'h6,8'h6,8'h6,8'h6,8'h22,8'h1a,8'h1a,8'h2b,8'h1a,8'h1a,8'h1a,8'h2b,8'h1a,8'h1a,8'h1a,8'h1a,8'h1a,8'h2b,8'h1a,8'h1a,8'h1a,8'h1a,8'h1a,8'h2b,8'h1a,8'h1a,8'h1a,8'h1a,8'h1a,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h1a,8'h21,8'h6,8'h2a,8'h1a,8'h1a,8'h21,8'h6,8'h6,8'h21,8'h1a,8'h1a,8'h1a,8'h1a,8'h1a,8'h1a,8'h1a,8'h1a,8'h1a,8'h1a,8'h1a,8'h21,8'h6,8'h2a,8'h1a,8'h2b,8'h1a,8'h1a,8'h2b,8'h1a,8'h1a,8'h1a,8'h2b,8'h2b,8'h1a,8'h1a,8'h2b,8'h2b,8'h1a,8'h1a,8'h1a,8'h1a,8'h1a,8'h1a,8'h1a,8'h1a,8'h2b,8'h1a,8'h1a,8'h1a,8'h1a,8'h1a,8'h1a,8'h2b,8'h1a,8'h1a,8'h1a,8'h1a,8'h1a,8'h1a,8'h1a,8'h1a,8'h1a,8'h1a,8'h1a,8'h1a,8'h1a,8'h2b,8'h1a,8'h1a,8'h2b,8'h1a,8'h1a,8'h1a,8'h1a,8'h1a,8'h2b,8'h1a,8'h1a,8'h21,8'h6,8'h6,8'h3,8'h2b,8'h1a,8'h1b,8'h6,8'h1b,8'h16,8'h1a,8'h21,8'h6,8'h6,8'h21,8'h2b,8'h1a,8'h9,8'h6,8'h6,8'h1b,8'h2b,8'h2b,8'h1a,8'h1a,8'h1a,8'h1a,8'h21,8'h22,8'h6,8'h6,8'h6,8'h6,8'h1b,8'h1a,8'h1a,8'h1a,8'h2b,8'h1a,8'h1a,8'h1a,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h18,8'h21,8'h6,8'h2a,8'h1a,8'h1a,8'h1a,8'h3,8'h6,8'h2a,8'h1a,8'h1a,8'h1a,8'h16,8'h1a,8'h1a,8'h1a,8'h16,8'h1a,8'h1a,8'h1a,8'h21,8'h6,8'h2a,8'h1a,8'h1a,8'h1a,8'h1a,8'h2b,8'h1a,8'h1a,8'h1a,8'h1a,8'h1a,8'h1a,8'h2b,8'h1a,8'h2b,8'h1a,8'h1a,8'h1a,8'h1a,8'h1a,8'h1a,8'h1a,8'h1a,8'h2b,8'h1a,8'h1a,8'h1a,8'h1a,8'h1a,8'h2b,8'h1a,8'h1a,8'h1a,8'h1a,8'h1a,8'h1a,8'h1a,8'h1a,8'h1a,8'h1a,8'h2b,8'h1a,8'h1a,8'h2b,8'h2b,8'h1a,8'h1a,8'h1a,8'h1a,8'h1a,8'h1a,8'h1a,8'h1a,8'h2b,8'h1a,8'h16,8'h7,8'h6,8'h21,8'h1a,8'h2b,8'h1a,8'h1a,8'h1a,8'h1a,8'h1a,8'h16,8'h6,8'h6,8'h21,8'h1a,8'h1a,8'h2b,8'h1a,8'ha,8'h6,8'h22,8'h1a,8'h2b,8'h1a,8'h1a,8'h1a,8'h1a,8'h21,8'h3,8'h1a,8'h1a,8'h3,8'h6,8'h2a,8'h1a,8'h1a,8'h1a,8'h1a,8'h1a,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h18,8'h21,8'h6,8'h2a,8'h1a,8'h18,8'h1a,8'h21,8'h6,8'h6,8'h1a,8'h1a,8'h1b,8'h6,8'h6,8'h6,8'h6,8'h9,8'h1a,8'h1a,8'h1a,8'h21,8'h6,8'h2a,8'h1a,8'h1b,8'h6,8'h6,8'h6,8'h1a,8'h1a,8'h18,8'h22,8'h6,8'h6,8'h6,8'h6,8'h21,8'h1a,8'h1a,8'ha,8'h6,8'h6,8'h6,8'h6,8'h6,8'h6,8'h6,8'h6,8'h6,8'h6,8'h3,8'h2b,8'h2b,8'h1a,8'h16,8'h6,8'h6,8'h6,8'h6,8'h22,8'h1b,8'h1a,8'h1a,8'h21,8'h6,8'h6,8'h6,8'h6,8'h6,8'h2,8'h1a,8'h1a,8'h1a,8'h1a,8'h1a,8'h2b,8'h1a,8'ha,8'h6,8'h2a,8'h1a,8'h1a,8'h1a,8'h1a,8'h1a,8'h1a,8'h1a,8'h18,8'ha,8'h6,8'h6,8'h1a,8'h1a,8'h1a,8'h1a,8'h1a,8'h1a,8'h6,8'h6,8'h21,8'h1a,8'h1a,8'h1a,8'h2b,8'h1a,8'h2b,8'h1a,8'h1a,8'h1a,8'h1b,8'h6,8'h6,8'h1b,8'h1a,8'h1a,8'h1a,8'h1a,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h18,8'h21,8'h6,8'h2a,8'h1a,8'h1a,8'h1a,8'h3,8'h6,8'h2a,8'h16,8'h1b,8'h6,8'h6,8'h21,8'h1a,8'h4,8'h6,8'h6,8'h16,8'h1a,8'h21,8'h6,8'h2a,8'h21,8'h6,8'h6,8'h3,8'h2b,8'h1a,8'h16,8'h7,8'h6,8'h21,8'h1a,8'h21,8'h6,8'h22,8'h1b,8'h1a,8'ha,8'h6,8'h2a,8'h1a,8'h16,8'h6,8'h6,8'h21,8'h1a,8'h1b,8'h6,8'h6,8'h1b,8'h2b,8'h21,8'h6,8'h6,8'h21,8'h1a,8'h3,8'h6,8'h22,8'h1a,8'h1a,8'h21,8'h6,8'h9,8'h1a,8'h1a,8'h9,8'h6,8'h2a,8'h1a,8'h1a,8'h1a,8'h1a,8'h2b,8'h1a,8'h9,8'h6,8'h2a,8'h1a,8'h1a,8'h1a,8'h1a,8'h1a,8'h1a,8'h1a,8'h1a,8'h9,8'h6,8'h2a,8'h1a,8'h1a,8'h1a,8'h1a,8'h1a,8'h1a,8'h22,8'h6,8'h21,8'h1a,8'h1a,8'h1a,8'h1a,8'h2b,8'h2b,8'h1a,8'h1a,8'h1a,8'h21,8'h6,8'h6,8'h1b,8'h1a,8'h1a,8'h1a,8'h1a,8'h1a,8'h1a,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h18,8'h21,8'h6,8'h2a,8'h16,8'h1a,8'h21,8'h6,8'h6,8'h21,8'h1a,8'h9,8'h6,8'h2a,8'h1a,8'h1a,8'h1a,8'h22,8'h6,8'h21,8'h1a,8'h21,8'h6,8'h6,8'h6,8'h6,8'h1b,8'h1a,8'h1a,8'h1a,8'ha,8'h6,8'h2a,8'h1a,8'h1a,8'h1a,8'h9,8'h6,8'h21,8'h1a,8'ha,8'h6,8'h2a,8'h1a,8'h1a,8'h9,8'h6,8'h2a,8'h1a,8'h1a,8'h6,8'h6,8'h3,8'h1a,8'h9,8'h6,8'h9,8'h1a,8'h1a,8'h1a,8'h22,8'h6,8'h21,8'h1a,8'h21,8'h6,8'h22,8'h1a,8'h1a,8'h1b,8'h6,8'h6,8'h1b,8'h1a,8'h1a,8'h1a,8'h1a,8'h1a,8'h17,8'h6,8'h2a,8'h1a,8'h1a,8'h1a,8'h1a,8'h1a,8'h1a,8'h1a,8'h18,8'hb,8'h6,8'h2a,8'h1a,8'h1a,8'h1a,8'h1a,8'h1a,8'h1a,8'h22,8'h6,8'h2,8'h1a,8'h1a,8'h2b,8'h2b,8'h1a,8'h1a,8'h1a,8'h1a,8'h1a,8'h6,8'h6,8'h2a,8'h1a,8'h1a,8'h1a,8'h1a,8'h1a,8'h2b,8'h1a,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h1a,8'h21,8'h6,8'h6,8'h6,8'h6,8'h6,8'h6,8'h1b,8'h1a,8'h1a,8'h6,8'h6,8'h21,8'h1a,8'h1a,8'h1a,8'h3,8'h6,8'h9,8'h1a,8'h21,8'h6,8'h6,8'h6,8'h2,8'h1a,8'h1a,8'h1a,8'h16,8'h6,8'h6,8'h6,8'h6,8'h6,8'h6,8'h6,8'h6,8'h2a,8'h1a,8'ha,8'h6,8'h2a,8'h1a,8'h1a,8'h3,8'h6,8'h2a,8'h1a,8'h1a,8'h9,8'h6,8'h21,8'h1a,8'h22,8'h6,8'h21,8'h1a,8'h1a,8'h1a,8'h21,8'h6,8'h2a,8'h1a,8'h21,8'h6,8'h22,8'h1a,8'h1a,8'h16,8'h6,8'h6,8'h1b,8'h1a,8'h1a,8'h1a,8'h2b,8'h1a,8'h9,8'h6,8'h2a,8'h1a,8'h1a,8'h1a,8'h1a,8'h9,8'h6,8'h3,8'h1a,8'h9,8'h6,8'h2,8'h1a,8'h1a,8'h1a,8'h2b,8'h1a,8'h1a,8'h6,8'h6,8'h21,8'h1a,8'h1a,8'h1a,8'h1a,8'h2b,8'h2b,8'h1a,8'h21,8'h6,8'h6,8'h6,8'h1a,8'h1a,8'h1a,8'h1a,8'h1a,8'h1a,8'h1a,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h1a,8'h21,8'h6,8'h22,8'h1a,8'h1a,8'h2b,8'h1a,8'h1a,8'h1a,8'h16,8'h22,8'h6,8'h21,8'h1a,8'h1a,8'h1a,8'h21,8'h6,8'h2,8'h1a,8'h21,8'h6,8'h6,8'h6,8'h6,8'h2,8'h1a,8'h1a,8'h1a,8'h6,8'h6,8'h3,8'h1a,8'h1a,8'h2b,8'h2b,8'h1a,8'h1a,8'h1a,8'h4,8'h6,8'h2a,8'h1a,8'h1a,8'h3,8'h6,8'h2a,8'h1a,8'h1a,8'h9,8'h6,8'h3,8'h1a,8'h22,8'h6,8'h21,8'h1a,8'h1a,8'h1a,8'h3,8'h6,8'h2a,8'h1a,8'h21,8'h6,8'h22,8'h2b,8'h1a,8'h16,8'h6,8'h6,8'h1b,8'h1a,8'h1a,8'h1a,8'h1a,8'h1a,8'ha,8'h6,8'h2a,8'h1a,8'h1a,8'h1a,8'h1a,8'h9,8'h6,8'h21,8'h1a,8'ha,8'h6,8'h6,8'h1a,8'h1a,8'h1a,8'h2b,8'h1a,8'h16,8'h6,8'h6,8'h21,8'h2b,8'h1a,8'h1a,8'h1a,8'h2b,8'h1a,8'h9,8'h6,8'h6,8'h1b,8'h1a,8'h1a,8'h1a,8'h1a,8'h1a,8'h1a,8'h2b,8'h2b,8'h1a,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h1a,8'h21,8'h6,8'h22,8'h1a,8'h1a,8'h1a,8'h2b,8'h1a,8'h1a,8'h1a,8'h9,8'h6,8'h3,8'h1a,8'h1a,8'h1a,8'h6,8'h6,8'h21,8'h1a,8'h21,8'h6,8'h2a,8'h2,8'h6,8'h6,8'h2,8'h1a,8'h1a,8'h3,8'h6,8'h2a,8'h1a,8'h1a,8'h2b,8'h1a,8'h1a,8'h1a,8'h1a,8'hb,8'h6,8'h2a,8'h1a,8'h1a,8'h4,8'h6,8'h2a,8'h1a,8'h1a,8'h9,8'h6,8'h21,8'h1a,8'h9,8'h6,8'h9,8'h2b,8'h1a,8'h1a,8'h6,8'h6,8'h3,8'h1a,8'h21,8'h6,8'h9,8'h1a,8'h1a,8'h1a,8'h6,8'h6,8'h1b,8'h1a,8'h1a,8'h1a,8'h1a,8'h1a,8'h21,8'h6,8'h6,8'h21,8'h1a,8'h1a,8'h1a,8'h9,8'h6,8'h21,8'h1a,8'h16,8'h6,8'h6,8'h2,8'h1a,8'h2b,8'h1a,8'h1a,8'h3,8'h6,8'h9,8'h1a,8'h1a,8'h1a,8'h1a,8'h1a,8'h1a,8'h16,8'h6,8'h6,8'h1b,8'h1a,8'h1a,8'h1a,8'h1a,8'h1a,8'h1a,8'h2b,8'h1a,8'h1a,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h1a,8'h21,8'h6,8'h2a,8'h1a,8'h1a,8'h1a,8'h2b,8'h1a,8'h1a,8'h1a,8'h1b,8'h6,8'h6,8'h21,8'h1a,8'h21,8'h6,8'h6,8'h1a,8'h16,8'h21,8'h6,8'h22,8'h1a,8'h3,8'h6,8'h6,8'h3,8'h1a,8'h1a,8'h6,8'h6,8'h2a,8'h2b,8'h1a,8'h2b,8'h2b,8'h1a,8'h1a,8'h4,8'h6,8'h2a,8'h1a,8'h1a,8'h3,8'h6,8'h2a,8'h1a,8'h1a,8'h9,8'h6,8'h3,8'h1a,8'h21,8'h6,8'h6,8'h21,8'h1a,8'h3,8'h6,8'h6,8'h1a,8'h1a,8'h21,8'h6,8'h22,8'h1a,8'h1a,8'h16,8'h6,8'h6,8'h1b,8'h1a,8'h2b,8'h1a,8'h1a,8'h1a,8'h1a,8'h4,8'h6,8'h6,8'h21,8'h1a,8'h1a,8'h9,8'h6,8'h3,8'h1a,8'h1a,8'h21,8'h22,8'h6,8'h3,8'h1a,8'h1a,8'h9,8'h6,8'h6,8'h1b,8'h2b,8'h2b,8'h1a,8'h1a,8'h1a,8'h1a,8'h9,8'h6,8'h22,8'h1a,8'h2b,8'h1a,8'h1a,8'h1a,8'h2b,8'h1a,8'h1a,8'h2b,8'h2b,8'h1a,8'h1a,8'h1a,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h1a,8'h21,8'h6,8'h22,8'h1a,8'h2b,8'h1a,8'h2b,8'h1a,8'h1a,8'h1a,8'h1a,8'h16,8'h6,8'h6,8'h6,8'h6,8'h6,8'h1a,8'h1a,8'h1a,8'h21,8'h6,8'h9,8'h1a,8'h1a,8'h9,8'h6,8'h6,8'h21,8'h1a,8'h1a,8'h6,8'h6,8'h6,8'h6,8'h6,8'h6,8'h1a,8'h1a,8'ha,8'h6,8'h9,8'h1a,8'h1a,8'h3,8'h6,8'h2a,8'h1a,8'h1a,8'h9,8'h6,8'h21,8'h1a,8'h1a,8'h1a,8'h22,8'h6,8'h6,8'h6,8'h22,8'h1b,8'h1a,8'h1a,8'h21,8'h6,8'h22,8'h1a,8'h1a,8'h16,8'h6,8'h6,8'h1b,8'h1a,8'h1a,8'h2b,8'h1a,8'h1a,8'h1a,8'h1a,8'h16,8'h6,8'h6,8'h6,8'h6,8'h6,8'h6,8'h3,8'h1a,8'h1a,8'h1a,8'h1a,8'h6,8'h6,8'h6,8'h6,8'h6,8'h9,8'h1a,8'h1a,8'h1a,8'h1a,8'h2b,8'h1a,8'h2b,8'h1a,8'h9,8'h6,8'h6,8'h6,8'h6,8'h6,8'h6,8'h3,8'h2b,8'h2b,8'h1a,8'h2b,8'h1a,8'h1a,8'h1a,8'h1a,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h1a,8'h1a,8'h1a,8'h1a,8'h1a,8'h1a,8'h2b,8'h2b,8'h1b,8'h1a,8'h1a,8'h1a,8'h1a,8'h1a,8'h2b,8'h1a,8'h1a,8'h2b,8'h1a,8'h1a,8'h1a,8'h1a,8'h1a,8'h1a,8'h1a,8'h2b,8'h1a,8'h1a,8'h1a,8'h1a,8'h1a,8'h1a,8'h1a,8'h1a,8'h1a,8'h1a,8'h1a,8'h1a,8'h1a,8'h1a,8'h1a,8'h2b,8'h1a,8'h1a,8'h1a,8'h2b,8'h1a,8'h1a,8'h1a,8'h1a,8'h1a,8'h1a,8'h2b,8'h1a,8'h1a,8'h1a,8'h1a,8'h1a,8'h1a,8'h1a,8'h1a,8'h1a,8'h1a,8'h1a,8'h1a,8'h1a,8'h1a,8'h1a,8'h1a,8'h1a,8'h1a,8'h2b,8'h1a,8'h1a,8'h1a,8'h2b,8'h1a,8'h1a,8'h1a,8'h1a,8'h2b,8'h1a,8'h1a,8'h1a,8'h1a,8'h2b,8'h1a,8'h1a,8'h1a,8'h1a,8'h1a,8'h1a,8'h1a,8'h1a,8'h1a,8'h1a,8'h1a,8'h1a,8'h2b,8'h2b,8'h1a,8'h1a,8'h2b,8'h1a,8'h1a,8'h1a,8'h1a,8'h1a,8'h1a,8'h1a,8'h1a,8'h1a,8'h2b,8'h1a,8'h1a,8'h1a,8'h1a,8'h1a,8'h1a,8'h1a,8'h1a,8'h1a,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h1a,8'h1a,8'h1a,8'h1a,8'h1a,8'h1a,8'h2b,8'h1a,8'h1a,8'h1a,8'h2b,8'h1a,8'h1a,8'h1a,8'h1a,8'h1a,8'h2b,8'h1a,8'h1a,8'h1a,8'h1a,8'h1a,8'h1a,8'h1a,8'h1a,8'h1a,8'h1a,8'h1a,8'h1a,8'h2b,8'h1a,8'h1a,8'h1a,8'h1a,8'h1a,8'h1a,8'h1a,8'h1a,8'h1a,8'h1a,8'h1a,8'h2b,8'h1a,8'h1a,8'h1a,8'h1a,8'h1a,8'h1a,8'h1a,8'h1a,8'h1a,8'h1a,8'h1a,8'h2b,8'h1a,8'h1a,8'h1a,8'h2b,8'h1a,8'h1a,8'h1a,8'h1a,8'h1a,8'h2b,8'h1a,8'h1a,8'h1a,8'h1a,8'h1a,8'h1a,8'h1a,8'h2b,8'h1a,8'h2b,8'h2b,8'h2b,8'h1a,8'h1a,8'h1a,8'h1a,8'h1a,8'h1a,8'h18,8'h1a,8'h2b,8'h1a,8'h1a,8'h1a,8'h1a,8'h1a,8'h1a,8'h1a,8'h1a,8'h1a,8'h1a,8'h1a,8'h1a,8'h1a,8'h1a,8'h1a,8'h1a,8'h1a,8'h1a,8'h1a,8'h1a,8'h1a,8'h1a,8'h2b,8'h1a,8'h1a,8'h1a,8'h1a,8'h1a,8'h1a,8'h2b,8'h1a,8'h1a,8'h1a,8'h1a,8'h1a,8'h1a,8'h1a,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h1a,8'h2b,8'h2b,8'h1a,8'h1a,8'h1a,8'h2b,8'h1a,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h1a,8'h1a,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h1a,8'h2b,8'h2b,8'h2b,8'h1a,8'h1a,8'h1a,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h1a,8'h1a,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h1a,8'h1a,8'h2b,8'h2b,8'h1a,8'h1a,8'h1a,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h1a,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h1a,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h1a,8'h1a,8'h1a,8'h1a,8'h1a,8'h1a,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h1a,8'h2b,8'h2b,8'h21,8'h6,8'h9,8'h1a,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h1a,8'h1a,8'h1a,8'h1a,8'h2b,8'h2b,8'h2b,8'h1a,8'h1a,8'h21,8'h6,8'h6,8'h6,8'h6,8'h6,8'h6,8'h1b,8'h1a,8'h1a,8'h21,8'h6,8'h22,8'h1a,8'h1a,8'h1a,8'h1a,8'h1a,8'h1a,8'h1a,8'h2b,8'h1a,8'h1a,8'h1a,8'h1a,8'h1a,8'h1a,8'h1a,8'h1a,8'h1a,8'h1a,8'h1a,8'h1a,8'h1a,8'h1a,8'h1a,8'h1a,8'h1a,8'h2b,8'h1a,8'h1a,8'h2b,8'h1a,8'h1a,8'h1a,8'h1a,8'h1a,8'h2b,8'h1a,8'h1a,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h1a,8'h1a,8'h1a,8'h1a,8'h1a,8'h1a,8'h1e,8'h1d,8'h1d,8'h11,8'ha,8'ha,8'ha,8'h1f,8'h1a,8'h1a,8'h1a,8'h1a,8'h1a,8'h16,8'h16,8'h1a,8'h2b,8'h1a,8'h1a,8'h1a,8'h2b,8'h1a,8'h1a,8'h1a,8'h1a,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h1a,8'h1a,8'h1b,8'h28,8'h2a,8'h28,8'h2a,8'h2a,8'h2a,8'h1a,8'h1a,8'h1a,8'h2b,8'h1a,8'h1a,8'h1a,8'h1a,8'h1a,8'h1a,8'h1a,8'h1a,8'h1a,8'h1a,8'h1a,8'h1a,8'h1a,8'h1a,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h1a,8'h1a,8'h1a,8'h1a,8'h2b,8'h2b,8'h2b,8'h1a,8'h1a,8'h21,8'h6,8'h9,8'h1a,8'h1a,8'h21,8'h6,8'h6,8'h21,8'h1a,8'h21,8'h6,8'h2a,8'h1a,8'h1a,8'h1a,8'h1a,8'h1a,8'h2b,8'h1a,8'h1a,8'h1a,8'h1a,8'h1a,8'h1a,8'h1a,8'h2b,8'h1a,8'h1a,8'h1a,8'h2b,8'h1a,8'h1a,8'h1a,8'h1a,8'h1a,8'h1a,8'h1a,8'h2b,8'h1a,8'h1a,8'h1a,8'h2b,8'h1a,8'h1a,8'h1a,8'h2b,8'h2b,8'h1a,8'h1a,8'h1a,8'h1a,8'h1a,8'h1a,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h1a,8'h1a,8'h1a,8'h1a,8'h1a,8'h1a,8'h1e,8'h1d,8'h1e,8'h1a,8'h16,8'h1e,8'ha,8'ha,8'h1f,8'h1a,8'h1a,8'h1a,8'h1a,8'h1e,8'h11,8'h21,8'h1a,8'h1a,8'h1a,8'h1a,8'h2b,8'h1a,8'h1a,8'h1a,8'h1a,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h1a,8'h2b,8'h1b,8'h2a,8'h28,8'h1a,8'h1a,8'h1b,8'h28,8'h2a,8'h27,8'h1a,8'h1a,8'h3,8'h2,8'h2a,8'h28,8'h2a,8'h1a,8'h1a,8'h1a,8'h1a,8'h1a,8'h1a,8'h1a,8'h1a,8'h1a,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h1a,8'h1a,8'h1a,8'h1a,8'h2b,8'h2b,8'h2b,8'h1a,8'h1a,8'h21,8'h6,8'h22,8'h1a,8'h1a,8'h1a,8'h3,8'h6,8'h6,8'h1b,8'h21,8'h6,8'h22,8'h1a,8'h1a,8'h1a,8'h1a,8'h1a,8'h2b,8'h1a,8'h1a,8'h1a,8'h1a,8'h1a,8'h1a,8'h1a,8'h1a,8'h2b,8'h1a,8'h1a,8'h1a,8'h1a,8'h1a,8'h2b,8'h1a,8'h1a,8'h2b,8'h1a,8'h1a,8'h2b,8'h1a,8'h1a,8'h2b,8'h1a,8'h1a,8'h1a,8'h2b,8'h1a,8'h1a,8'h1a,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h1a,8'h1a,8'h2b,8'h1a,8'h1a,8'h1a,8'h1a,8'h1e,8'h1d,8'h1e,8'h18,8'h1a,8'h1a,8'h1e,8'h1e,8'h1e,8'h1a,8'h1a,8'h1a,8'h1e,8'ha,8'ha,8'h1b,8'h1a,8'h1a,8'h1a,8'h2b,8'h2b,8'h1a,8'h1a,8'h2b,8'h1a,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h1a,8'h1a,8'h1b,8'h28,8'h27,8'h1a,8'h1a,8'h1a,8'h27,8'h2a,8'h27,8'h1a,8'h21,8'h21,8'h1a,8'h1a,8'h27,8'h28,8'h2a,8'h1a,8'h1a,8'h1a,8'h1a,8'h1a,8'h1a,8'h1a,8'h1a,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h1a,8'h1a,8'h1a,8'h1a,8'h2b,8'h2b,8'h2b,8'h1a,8'h1a,8'h21,8'h6,8'h22,8'h1a,8'h1a,8'h1a,8'h21,8'h6,8'h6,8'h1a,8'h1,8'h6,8'h2a,8'h1a,8'h1a,8'h21,8'h6,8'h22,8'h6,8'h6,8'h6,8'h1b,8'h1a,8'h21,8'h6,8'h22,8'h1a,8'h1a,8'h16,8'h6,8'h6,8'h21,8'h1a,8'h1a,8'h6,8'h6,8'h6,8'h6,8'h6,8'h1b,8'h1a,8'h2b,8'h21,8'h6,8'h6,8'h6,8'h6,8'h6,8'h21,8'h1a,8'h1a,8'h2b,8'h2b,8'h1a,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h1a,8'h1a,8'h2b,8'h1a,8'h1a,8'h1a,8'h1a,8'h1f,8'h1d,8'h1e,8'h1a,8'h1a,8'h1a,8'h1f,8'h1d,8'h1d,8'h1a,8'h1a,8'h21,8'ha,8'h1d,8'ha,8'h21,8'h1a,8'h1a,8'h1a,8'h2b,8'h2b,8'h1a,8'h1a,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h1a,8'h2b,8'h1b,8'h2a,8'h28,8'h1a,8'h1a,8'h1a,8'h1b,8'h2a,8'h2a,8'h1a,8'h1a,8'h1a,8'h1a,8'h1a,8'h1a,8'h2a,8'h2a,8'h1b,8'h1a,8'h1a,8'h1a,8'h1a,8'h1a,8'h1a,8'h1a,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h1a,8'h1a,8'h1a,8'h1a,8'h2b,8'h2b,8'h2b,8'h1a,8'h1a,8'h21,8'h6,8'h22,8'h1a,8'h1a,8'h1a,8'h3,8'h6,8'h6,8'h1a,8'h21,8'h6,8'h2a,8'h1a,8'h1a,8'h1a,8'h1a,8'h1a,8'h1a,8'h3,8'h6,8'h6,8'h1a,8'h1b,8'h6,8'h6,8'h1a,8'h1a,8'h1b,8'h6,8'h6,8'h1a,8'h16,8'h6,8'h6,8'h21,8'h2b,8'h21,8'h6,8'h6,8'h1b,8'h2b,8'h21,8'h6,8'h6,8'h1a,8'h1a,8'h1a,8'h1a,8'h1a,8'h1a,8'h1a,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h1a,8'h2b,8'h1a,8'h1a,8'h1a,8'h1a,8'h1f,8'ha,8'h1e,8'h1a,8'h1a,8'h1a,8'h1e,8'ha,8'h1e,8'h1a,8'h21,8'ha,8'h1e,8'h1e,8'h1d,8'h21,8'h1a,8'h1a,8'h1a,8'h2b,8'h2b,8'h1a,8'h1a,8'h2b,8'h1a,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h1a,8'h1b,8'h28,8'h28,8'h1a,8'h1a,8'h1a,8'h1b,8'h28,8'h2a,8'h1a,8'h1a,8'h1a,8'h1a,8'h1a,8'h1b,8'h2a,8'h2a,8'h1b,8'h1a,8'h2b,8'h1a,8'h1a,8'h1a,8'h1a,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h1a,8'h1a,8'h1a,8'h1a,8'h2b,8'h2b,8'h2b,8'h1a,8'h1a,8'h21,8'h6,8'h2a,8'h1a,8'h1a,8'h21,8'h6,8'h6,8'h3,8'h1a,8'h1,8'h6,8'h2a,8'h1a,8'h1a,8'h1a,8'h1a,8'h1a,8'h1a,8'h1a,8'h6,8'h6,8'h1b,8'h1a,8'h17,8'h6,8'h2,8'h1a,8'h3,8'h6,8'h2a,8'h1a,8'hb,8'h6,8'h2a,8'h1a,8'h2b,8'h1a,8'h9,8'h6,8'h3,8'h1a,8'h21,8'h6,8'h6,8'h1a,8'h1a,8'h1a,8'h1a,8'h1a,8'h1a,8'h1a,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h1a,8'h1a,8'h2b,8'h1a,8'h1a,8'h1a,8'h1a,8'h1f,8'ha,8'h1e,8'h1a,8'h16,8'h1f,8'ha,8'ha,8'h1f,8'h1a,8'h1a,8'h1a,8'h16,8'h1e,8'h1d,8'h1e,8'h1a,8'h1a,8'h1a,8'h1a,8'h2b,8'h1a,8'h1a,8'h1a,8'h1a,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h1b,8'h2a,8'h27,8'h1a,8'h1a,8'h1b,8'h2a,8'h2a,8'h21,8'h1a,8'h1a,8'h1a,8'h1a,8'h1a,8'h28,8'h2a,8'h21,8'h1a,8'h1a,8'h2b,8'h1a,8'h1a,8'h1a,8'h1a,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h1a,8'h1a,8'h1a,8'h1a,8'h2b,8'h2b,8'h2b,8'h1a,8'h1a,8'h21,8'h6,8'h6,8'h6,8'h6,8'h6,8'h6,8'h1b,8'h1a,8'h1a,8'h21,8'h6,8'h6,8'h1a,8'h1a,8'h1a,8'h22,8'h6,8'h6,8'h6,8'h6,8'h6,8'h1b,8'h1a,8'ha,8'h6,8'h22,8'h1a,8'h9,8'h6,8'h3,8'h1a,8'h9,8'h6,8'h6,8'h6,8'h6,8'h6,8'h6,8'h6,8'h2,8'h1a,8'h21,8'h6,8'h6,8'h1a,8'h1a,8'h1a,8'h1a,8'h1a,8'h1a,8'h1a,8'h2b,8'h1a,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h1a,8'h1a,8'h2b,8'h1a,8'h1a,8'h1a,8'h1a,8'h1f,8'ha,8'h1d,8'h11,8'ha,8'ha,8'ha,8'h16,8'h1a,8'h1a,8'h1a,8'h1a,8'h1a,8'h1e,8'h1d,8'h1e,8'h1a,8'h1a,8'h1a,8'h1a,8'h2b,8'h1a,8'h1a,8'h1a,8'h1a,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h1a,8'h1a,8'h1b,8'h2a,8'h2a,8'h28,8'h2a,8'h2a,8'h2a,8'h1b,8'h1a,8'h1a,8'h2b,8'h1a,8'h1a,8'h2a,8'h2a,8'h2a,8'h1a,8'h1a,8'h1a,8'h1a,8'h1a,8'h1a,8'h1a,8'h1a,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h1a,8'h1a,8'h1a,8'h2b,8'h2b,8'h2b,8'h1a,8'h1a,8'h21,8'h6,8'h9,8'h1a,8'h1a,8'h1a,8'h1a,8'h2b,8'h1a,8'h1a,8'h21,8'h6,8'h2a,8'h1a,8'h1a,8'h22,8'h6,8'h9,8'h1a,8'h16,8'h6,8'h6,8'h1b,8'h1a,8'h16,8'h6,8'h6,8'h6,8'h6,8'h6,8'h1b,8'h1a,8'h6,8'h6,8'h3,8'h1a,8'h1a,8'h1a,8'h1a,8'h2b,8'h1a,8'h2b,8'h21,8'h6,8'h6,8'h1a,8'h1a,8'h1a,8'h1a,8'h1a,8'h1a,8'h1a,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h1a,8'h1a,8'h2b,8'h1a,8'h1a,8'h1a,8'h1a,8'h1f,8'ha,8'h1e,8'h1a,8'h1a,8'h1a,8'h1a,8'h1a,8'h1a,8'h1a,8'h1a,8'h1a,8'h1a,8'h1d,8'h1d,8'h1f,8'h1a,8'h1a,8'h1a,8'h2b,8'h2b,8'h1a,8'h1a,8'h1a,8'h1a,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h1a,8'h2b,8'h1b,8'h2a,8'h28,8'h1a,8'h1a,8'h1a,8'h1a,8'h2b,8'h1a,8'h1a,8'h2b,8'h21,8'h2a,8'h28,8'h1a,8'h1a,8'h1a,8'h1a,8'h1a,8'h2b,8'h2b,8'h1a,8'h1a,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h1a,8'h1a,8'h1a,8'h2b,8'h2b,8'h2b,8'h1a,8'h1a,8'h21,8'h6,8'h2a,8'h1a,8'h1a,8'h1a,8'h1a,8'h2b,8'h2b,8'h1a,8'h21,8'h6,8'h22,8'h1a,8'h16,8'h6,8'h6,8'h1b,8'h1a,8'h16,8'h6,8'h6,8'h1b,8'h1a,8'h1a,8'h9,8'h6,8'h6,8'h6,8'h9,8'h1a,8'h2b,8'ha,8'h6,8'h2a,8'h1a,8'h1a,8'h1a,8'h1a,8'h1a,8'h1a,8'h2b,8'h21,8'h6,8'h6,8'h1a,8'h1a,8'h1a,8'h1a,8'h1a,8'h1a,8'h1a,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h1a,8'h1a,8'h1a,8'h1a,8'h1a,8'h1a,8'h1a,8'h1f,8'ha,8'h1e,8'h1a,8'h1a,8'h1a,8'h1a,8'h1a,8'h1a,8'h1a,8'h1a,8'h1a,8'h1a,8'h1e,8'h1d,8'h1e,8'h1a,8'h1a,8'h1a,8'h2b,8'h1a,8'h1a,8'h1a,8'h2b,8'h1a,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h1a,8'h2b,8'h1b,8'h2a,8'h27,8'h1a,8'h1a,8'h1a,8'h1a,8'h1a,8'h1a,8'h1a,8'h1b,8'h2a,8'h2a,8'h1a,8'h1a,8'h1a,8'h1a,8'h1a,8'h1a,8'h1a,8'h1a,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h1a,8'h1a,8'h1a,8'h2b,8'h2b,8'h2b,8'h1a,8'h1a,8'h21,8'h6,8'h9,8'h1a,8'h1a,8'h1a,8'h1a,8'h1a,8'h1a,8'h1a,8'h21,8'h6,8'h6,8'h1a,8'h1a,8'h22,8'h6,8'h21,8'h1a,8'h16,8'h6,8'h6,8'h1b,8'h1a,8'h1a,8'h1b,8'h6,8'h6,8'h6,8'h21,8'h2b,8'h1a,8'h16,8'h6,8'h6,8'h2a,8'h1a,8'h1a,8'h1a,8'h1a,8'h1a,8'h2b,8'h21,8'h6,8'h6,8'h1a,8'h1a,8'h1a,8'h1a,8'h1a,8'h1a,8'h1a,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h1a,8'h1a,8'h1a,8'h1a,8'h1a,8'h1a,8'h1a,8'h1f,8'ha,8'h1e,8'h1a,8'h1a,8'h1a,8'h1a,8'h1a,8'h1a,8'h1a,8'h1a,8'h1a,8'h1a,8'h12,8'ha,8'h21,8'h1a,8'h1a,8'h2b,8'h2b,8'h1a,8'h1a,8'h1a,8'h2b,8'h1a,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h1a,8'h2b,8'h1b,8'h2a,8'h28,8'h1a,8'h1a,8'h1a,8'h1a,8'h1a,8'h1a,8'h1a,8'h21,8'h2a,8'h21,8'h1a,8'h1a,8'h1a,8'h1a,8'h1a,8'h2b,8'h2b,8'h1a,8'h1a,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h1a,8'h1a,8'h1a,8'h2b,8'h2b,8'h2b,8'h1a,8'h1a,8'h21,8'h6,8'h2a,8'h1a,8'h1a,8'h1a,8'h2b,8'h1a,8'h1a,8'h1a,8'h1a,8'h3,8'h6,8'h6,8'h16,8'h16,8'h6,8'h6,8'h6,8'h6,8'h6,8'h6,8'h1b,8'h1a,8'h1a,8'h1a,8'h9,8'h6,8'h6,8'h1a,8'h1a,8'h1a,8'h2b,8'h1a,8'h6,8'h22,8'h6,8'h6,8'h6,8'h22,8'h1b,8'h2b,8'h21,8'h6,8'h6,8'h1a,8'h1a,8'h1a,8'h1a,8'h1a,8'h2b,8'h1a,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h1a,8'h2b,8'h1a,8'h1a,8'h1a,8'h1a,8'h1a,8'h1f,8'ha,8'ha,8'h1a,8'h1a,8'h1a,8'h1a,8'h1a,8'h1a,8'h1a,8'h1a,8'h1a,8'h1a,8'ha,8'ha,8'h21,8'h1a,8'h2b,8'h2b,8'h1a,8'h1a,8'h1a,8'h1a,8'h2b,8'h1a,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h1a,8'h2b,8'h1b,8'h2a,8'h28,8'h1a,8'h1a,8'h2b,8'h1a,8'h1a,8'h1a,8'h1a,8'h21,8'h2a,8'h2a,8'h2a,8'h2a,8'h2a,8'h2a,8'h21,8'h1a,8'h2b,8'h2b,8'h1a,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h1a,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h1a,8'h1a,8'h1a,8'h2b,8'h2b,8'h2b,8'h1a,8'h1a,8'h1a,8'h18,8'h1a,8'h1a,8'h1a,8'h1a,8'h2b,8'h2b,8'h1a,8'h1a,8'h1a,8'h2b,8'h1a,8'h1a,8'h2b,8'h2b,8'h2b,8'h1a,8'h1a,8'h1a,8'h1a,8'h1a,8'h1a,8'h1a,8'h1a,8'h1a,8'h3,8'h6,8'h2,8'h1a,8'h2b,8'h1a,8'h2b,8'h2b,8'h1a,8'h1a,8'h2b,8'h1a,8'h1a,8'h1a,8'h1a,8'h2b,8'h1a,8'h1a,8'h1a,8'h1a,8'h1a,8'h1a,8'h1a,8'h1a,8'h2b,8'h1a,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h1a,8'h1a,8'h1a,8'h1a,8'h1a,8'h1a,8'h1a,8'h1a,8'h1a,8'h1a,8'h2b,8'h1a,8'h1a,8'h1a,8'h2b,8'h2b,8'h1a,8'h1a,8'h16,8'h1a,8'h1a,8'h1a,8'h2b,8'h2b,8'h1a,8'h1a,8'h1a,8'h1a,8'h2b,8'h1a,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h1a,8'h1a,8'h1a,8'h1a,8'h1a,8'h1a,8'h1a,8'h1a,8'h1a,8'h1a,8'h1a,8'h1a,8'h1a,8'h1a,8'h1a,8'h1a,8'h1a,8'h1a,8'h1a,8'h2b,8'h2b,8'h1a,8'h1a,8'h1a,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h1a,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h1a,8'h1a,8'h1a,8'h2b,8'h2b,8'h2b,8'h1a,8'h1a,8'h1a,8'h1a,8'h1a,8'h1a,8'h1a,8'h1a,8'h1a,8'h1a,8'h1a,8'h1a,8'h1a,8'h2b,8'h2b,8'h2b,8'h1a,8'h1a,8'h1a,8'h1a,8'h1a,8'h1a,8'h1a,8'h1a,8'h1a,8'h1a,8'h1a,8'h1b,8'h6,8'h6,8'h1b,8'h1a,8'h2b,8'h1a,8'h1a,8'h1a,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h1a,8'h1a,8'h2b,8'h1a,8'h1a,8'h1a,8'h1a,8'h1a,8'h1a,8'h1a,8'h1a,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h1a,8'h2b,8'h1a,8'h1a,8'h1a,8'h1a,8'h1a,8'h1a,8'h1a,8'h1a,8'h1a,8'h1a,8'h1a,8'h2b,8'h2b,8'h2b,8'h1a,8'h1a,8'h1a,8'h1a,8'h1a,8'h1a,8'h1a,8'h2b,8'h2b,8'h2b,8'h1a,8'h1a,8'h1a,8'h1a,8'h2b,8'h1a,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h1a,8'h1a,8'h1a,8'h1a,8'h1a,8'h1a,8'h2b,8'h1a,8'h1a,8'h1a,8'h1a,8'h1a,8'h1a,8'h1a,8'h1a,8'h1a,8'h1a,8'h2b,8'h2b,8'h2b,8'h1a,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h1a,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h1a,8'h1a,8'h1a,8'h2b,8'h2b,8'h2b,8'h1a,8'h1a,8'h1a,8'h1a,8'h1a,8'h1a,8'h1a,8'h1a,8'h2b,8'h1a,8'h1a,8'h1a,8'h2b,8'h1a,8'h1a,8'h1a,8'h2b,8'h2b,8'h2b,8'h1a,8'h1a,8'h1a,8'h1a,8'h1a,8'h1a,8'h9,8'h6,8'h6,8'h6,8'h1b,8'h1a,8'h1a,8'h1a,8'h1a,8'h1a,8'h1a,8'h1a,8'h1a,8'h2b,8'h1a,8'h1a,8'h2b,8'h1a,8'h1a,8'h1a,8'h2b,8'h1a,8'h1a,8'h2b,8'h2b,8'h1a,8'h1a,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h1a,8'h2b,8'h1a,8'h1a,8'h1a,8'h1a,8'h1a,8'h1a,8'h1a,8'h1a,8'h1a,8'h1a,8'h2b,8'h1a,8'h1a,8'h1a,8'h1a,8'h2b,8'h1a,8'h1a,8'h1a,8'h1a,8'h1a,8'h1a,8'h1a,8'h2b,8'h1a,8'h1a,8'h1a,8'h1a,8'h2b,8'h1a,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h1a,8'h1a,8'h1a,8'h1a,8'h1a,8'h1a,8'h2b,8'h2b,8'h2b,8'h1a,8'h1a,8'h1a,8'h1a,8'h2b,8'h1a,8'h1a,8'h1a,8'h2b,8'h2b,8'h1a,8'h1a,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h1a,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h1a,8'h1a,8'h1a,8'h2b,8'h2b,8'h2b,8'h1a,8'h1a,8'h1a,8'h1a,8'h1a,8'h1a,8'h1a,8'h1a,8'h1a,8'h2b,8'h1a,8'h1a,8'h1a,8'h1a,8'h1a,8'h1a,8'h1a,8'h1a,8'h1a,8'h1a,8'h1a,8'h1a,8'h1a,8'h1a,8'h1a,8'h1a,8'h1a,8'h1a,8'h1a,8'h1a,8'h1a,8'h1a,8'h1a,8'h1a,8'h1a,8'h1a,8'h1a,8'h2b,8'h2b,8'h1a,8'h2b,8'h2b,8'h1a,8'h2b,8'h2b,8'h1a,8'h1a,8'h1a,8'h2b,8'h2b,8'h1a,8'h1a,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h1a,8'h1a,8'h1a,8'h1a,8'h1a,8'h1a,8'h1a,8'h1a,8'h1a,8'h1a,8'h1a,8'h1a,8'h1a,8'h1a,8'h1a,8'h1a,8'h1a,8'h1a,8'h1a,8'h1a,8'h1a,8'h1a,8'h1a,8'h1a,8'h1a,8'h1a,8'h1a,8'h1a,8'h1a,8'h1a,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h1a,8'h1a,8'h1a,8'h2b,8'h1a,8'h1a,8'h1a,8'h1a,8'h1a,8'h1a,8'h1a,8'h1a,8'h1a,8'h1a,8'h1a,8'h1a,8'h1a,8'h1a,8'h2b,8'h2b,8'h2b,8'h1a,8'h1a,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h1a,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h1a,8'h1a,8'h1a,8'h2b,8'h2b,8'h2b,8'h1a,8'h1a,8'h1a,8'h1a,8'h1a,8'h1a,8'h1a,8'h1a,8'h2b,8'h1a,8'h1a,8'h1a,8'h1a,8'h1a,8'h1a,8'h1a,8'h1a,8'h1a,8'h1a,8'h1a,8'h1a,8'h1a,8'h1a,8'h1a,8'h1a,8'h1a,8'h1a,8'h1a,8'h1a,8'h2b,8'h1a,8'h1a,8'h1a,8'h1a,8'h2b,8'h1a,8'h1a,8'h1a,8'h2b,8'h1a,8'h2b,8'h1a,8'h1a,8'h1a,8'h1a,8'h2b,8'h1a,8'h1a,8'h2b,8'h2b,8'h1a,8'h1a,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h1a,8'h1a,8'h1a,8'h1a,8'h1a,8'h1a,8'h1a,8'h1a,8'h1a,8'h1a,8'h1a,8'h1a,8'h1a,8'h1a,8'h1a,8'h1a,8'h1a,8'h1a,8'h1a,8'h1a,8'h1a,8'h1a,8'h1a,8'h1a,8'h1a,8'h1a,8'h1a,8'h1a,8'h1a,8'h1a,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h1a,8'h1a,8'h1a,8'h1a,8'h1a,8'h1a,8'h1a,8'h1a,8'h1a,8'h1a,8'h2b,8'h2b,8'h1a,8'h1a,8'h1a,8'h1a,8'h2b,8'h1a,8'h1a,8'h1a,8'h2b,8'h1a,8'h1a,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h1a,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h1a,8'h2b,8'h1a,8'h1a,8'h1a,8'h1a,8'h1a,8'h1a,8'h1a,8'h2b,8'h2b,8'h1a,8'h1a,8'h1a,8'h1a,8'h1a,8'h1a,8'h1a,8'h1a,8'h1a,8'h2b,8'h1a,8'h2b,8'h1a,8'h1a,8'h2b,8'h1a,8'h1a,8'h2b,8'h1a,8'h1a,8'h2b,8'h2b,8'h1a,8'h1a,8'h1a,8'h2b,8'h1a,8'h1a,8'h1a,8'h2b,8'h2b,8'h1a,8'h1a,8'h1a,8'h1a,8'h1a,8'h1a,8'h1a,8'h1a,8'h1a,8'h1a,8'h1a,8'h1a,8'h1a,8'h1a,8'h1a,8'h1a,8'h1a,8'h1a,8'h1a,8'h1a,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h1a,8'h1a,8'h1a,8'h1a,8'h1a,8'h1a,8'h2b,8'h1a,8'h1a,8'h1a,8'h1a,8'h2b,8'h2b,8'h1a,8'h2b,8'h2b,8'h1a,8'h1a,8'h1a,8'h1a,8'h1a,8'h1a,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h1a,8'h1a,8'h1a,8'h1a,8'h1a,8'h1a,8'h1a,8'h1a,8'h1a,8'h1a,8'h2b,8'h1a,8'h1a,8'h2b,8'h1a,8'h1a,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h1a,8'h1a,8'h1a,8'h1a,8'h1a,8'h1a,8'h1a,8'h1a,8'h1a,8'h2b,8'h1a,8'h1a,8'h1a,8'h1a,8'h1a,8'h1a,8'h1a,8'h1a,8'h2b,8'h1a,8'h2b,8'h1a,8'h1a,8'h1a,8'h1a,8'h1a,8'h1a,8'h1a,8'h1a,8'h2b,8'h1a,8'h2b,8'h1a,8'h16,8'h2b,8'h2b,8'h1a,8'h1a,8'h2b,8'h1a,8'h1a,8'h1a,8'h2b,8'h1a,8'h1a,8'h1a,8'h1a,8'h1a,8'h1a,8'h1a,8'h1a,8'h1a,8'h1a,8'h1a,8'h1a,8'h1a,8'h1a,8'h1a,8'h1a,8'h1a,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h1a,8'h1a,8'h1a,8'h1a,8'h1a,8'h1a,8'h2b,8'h1a,8'h1a,8'h2b,8'h1a,8'h1a,8'h2b,8'h1a,8'h1a,8'h1a,8'h2b,8'h1a,8'h1a,8'h1a,8'h1a,8'h1a,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h1a,8'h1a,8'h1a,8'h2b,8'h1a,8'h1a,8'h1a,8'h2b,8'h2b,8'h1a,8'h1a,8'h2b,8'h2b,8'h2b,8'h1a,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h1a,8'h1a,8'h1a,8'h1a,8'h1a,8'h1a,8'h1a,8'h2b,8'h2b,8'h1a,8'h1a,8'h1a,8'h1a,8'h1a,8'h1a,8'h1a,8'h1a,8'h1a,8'h2b,8'h2b,8'h2b,8'h2b,8'h1a,8'h2b,8'h1a,8'h1a,8'h1a,8'h1a,8'h1a,8'h1a,8'h2b,8'h1a,8'h1a,8'h1a,8'h1a,8'h1a,8'h2b,8'h1a,8'h1a,8'h2b,8'h2b,8'h2b,8'h1a,8'h1a,8'h1a,8'h2b,8'h1a,8'h1a,8'h1a,8'h2b,8'h1a,8'h2b,8'h1a,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h1a,8'h1a,8'h2b,8'h2b,8'h1a,8'h1a,8'h1a,8'h1a,8'h1a,8'h1a,8'h1a,8'h1a,8'h1a,8'h1a,8'h2b,8'h1a,8'h1a,8'h1a,8'h1a,8'h1a,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h1a,8'h1a,8'h1a,8'h1a,8'h1a,8'h1a,8'h1a,8'h1a,8'h1a,8'h1a,8'h1a,8'h1a,8'h1a,8'h2b,8'h1a,8'h1a,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h1a,8'h1a,8'h1a,8'h1a,8'h1a,8'h2b,8'h2,8'h6,8'h6,8'h6,8'h6,8'h6,8'h1b,8'h1a,8'h1a,8'h1a,8'h1a,8'h1a,8'h2b,8'h1a,8'h2b,8'h1a,8'h1a,8'h1a,8'h1a,8'h1a,8'h1a,8'h2b,8'h2b,8'h1a,8'h2b,8'h1a,8'h1a,8'h1a,8'h2b,8'h1a,8'h2b,8'h1a,8'h1a,8'h1a,8'h1a,8'h1a,8'h1a,8'h1a,8'h2b,8'h2b,8'h2b,8'h2b,8'h1a,8'h1a,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h1a,8'h2b,8'h1a,8'h1a,8'h1a,8'h1a,8'h1a,8'h1a,8'h3,8'h6,8'h22,8'h1a,8'h2b,8'h1a,8'h16,8'h6,8'h6,8'h21,8'h1a,8'h2b,8'h2b,8'h1a,8'h1a,8'h1a,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h1a,8'h1a,8'h1a,8'h21,8'h6,8'h6,8'h1b,8'h1a,8'h2b,8'h1a,8'h21,8'h6,8'h6,8'h1b,8'h1a,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h1a,8'h1a,8'h1a,8'h1a,8'h9,8'h6,8'h9,8'h1a,8'h1a,8'h1a,8'h21,8'h1b,8'h1a,8'h21,8'h6,8'h2a,8'h2b,8'h2b,8'h2b,8'h1a,8'h1a,8'h1a,8'h1a,8'h1a,8'h1a,8'h1a,8'h2b,8'h1a,8'h1a,8'h2b,8'h1a,8'h1a,8'h1a,8'h1a,8'h1a,8'h1a,8'h1a,8'h1a,8'h1a,8'h1a,8'h1a,8'h16,8'h2b,8'h2b,8'h1a,8'h1a,8'h2b,8'h2b,8'h1a,8'h1a,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h1a,8'h1a,8'h1a,8'h1a,8'h2b,8'h1a,8'h1a,8'h1a,8'h4,8'h6,8'h9,8'h1a,8'h1a,8'h1a,8'h1a,8'h7,8'h6,8'h21,8'h1a,8'h2b,8'h1a,8'h1a,8'h1a,8'h1a,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h1a,8'h1a,8'h21,8'h6,8'h6,8'h1a,8'h1a,8'h1a,8'h1a,8'h1b,8'h6,8'h6,8'h1b,8'h2b,8'h1a,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h1a,8'h1a,8'h1a,8'h1b,8'h22,8'h6,8'h21,8'h1a,8'h2b,8'h2b,8'h1a,8'h1a,8'h1a,8'h21,8'h6,8'h2a,8'h1a,8'h2b,8'h1a,8'h1a,8'h1a,8'h1a,8'h1a,8'h1a,8'h1a,8'h1a,8'h2b,8'h2b,8'h2b,8'h1a,8'h1a,8'h1a,8'h1a,8'h1a,8'h1a,8'h1a,8'h1a,8'h1a,8'h1a,8'h1a,8'h1a,8'h1a,8'h1a,8'h1a,8'h1a,8'h2b,8'h1a,8'h2b,8'h2b,8'h1a,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h1a,8'h1a,8'h1a,8'h1a,8'h2b,8'h1a,8'h1a,8'h1a,8'ha,8'h6,8'h22,8'h1a,8'h1a,8'h1a,8'h16,8'h6,8'h6,8'h21,8'h1a,8'h1a,8'h2b,8'h2b,8'h1a,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h1a,8'h1a,8'h21,8'h6,8'h6,8'h1a,8'h1a,8'h1a,8'h1a,8'h1b,8'h6,8'h6,8'h1b,8'h2b,8'h1a,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h1a,8'h1a,8'h6,8'h6,8'h9,8'h2b,8'h1a,8'h1a,8'h1a,8'h1a,8'h1a,8'h21,8'h6,8'h6,8'h22,8'h6,8'h6,8'h1b,8'h1a,8'h16,8'h6,8'h6,8'h6,8'h6,8'h9,8'h1a,8'h1a,8'h2b,8'h21,8'h6,8'h6,8'h6,8'h6,8'h6,8'h9,8'h1a,8'h1a,8'h1a,8'h1a,8'h1a,8'h22,8'h6,8'h6,8'h6,8'h22,8'h21,8'h1a,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h1a,8'h1a,8'h1a,8'h1a,8'h1a,8'h1a,8'h1a,8'h1a,8'ha,8'h6,8'h22,8'h1a,8'h1a,8'h1a,8'h16,8'h7,8'h6,8'h21,8'h1a,8'h1a,8'h2b,8'h2b,8'h1a,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h1a,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h1a,8'h1a,8'h21,8'h6,8'h6,8'h1a,8'h1a,8'h1a,8'h1a,8'h1b,8'h6,8'h6,8'h1b,8'h1a,8'h1a,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h1a,8'h1a,8'h21,8'h6,8'h6,8'h6,8'h6,8'h6,8'h1b,8'h1a,8'h1a,8'h21,8'h6,8'h2a,8'h1a,8'h1a,8'h2b,8'h1a,8'h1b,8'h6,8'h6,8'h21,8'h1a,8'h3,8'h6,8'h6,8'h1a,8'h1a,8'h4,8'h22,8'h22,8'h1a,8'h1a,8'h9,8'h6,8'h22,8'h1a,8'h1a,8'h16,8'h6,8'h6,8'h21,8'h1a,8'h21,8'h6,8'h22,8'h1b,8'h1a,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h1a,8'h1a,8'h1a,8'h1a,8'h1a,8'h2b,8'h1a,8'h1a,8'ha,8'h6,8'h22,8'h1a,8'h1a,8'h1a,8'h18,8'h6,8'h6,8'h21,8'h1a,8'h1a,8'h1a,8'h2b,8'h1a,8'h1a,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h1a,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h1a,8'h1a,8'h21,8'h6,8'h6,8'h1a,8'h1a,8'h1a,8'h1a,8'h1b,8'h6,8'h6,8'h1b,8'h1a,8'h1a,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h1a,8'h1a,8'h16,8'h6,8'h6,8'h6,8'h6,8'h6,8'h21,8'h1a,8'h21,8'h6,8'h2a,8'h1a,8'h1a,8'h2b,8'h1a,8'h9,8'h6,8'h2a,8'h1a,8'h1a,8'h1a,8'h22,8'h6,8'h21,8'h1a,8'h21,8'h6,8'h22,8'h1a,8'h1a,8'h1b,8'h6,8'h6,8'h1b,8'h1a,8'h3,8'h6,8'h9,8'h1a,8'h1a,8'h1a,8'h9,8'h6,8'h21,8'h1a,8'h1a,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h1a,8'h1a,8'h1a,8'h1a,8'h1a,8'h2b,8'h1a,8'h1a,8'ha,8'h6,8'h22,8'h1a,8'h1a,8'h1a,8'h18,8'h7,8'h6,8'h21,8'h1a,8'h1a,8'h1a,8'h2b,8'h1a,8'h1a,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h1a,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h1a,8'h18,8'h21,8'h6,8'h6,8'h6,8'h6,8'h6,8'h6,8'h6,8'h6,8'h2a,8'h1b,8'h1a,8'h1a,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h1a,8'h2b,8'h1a,8'h1a,8'h1a,8'h1a,8'h16,8'h22,8'h6,8'h6,8'h1a,8'h21,8'h6,8'h2a,8'h1a,8'h2b,8'h2b,8'h1a,8'h6,8'h6,8'h21,8'h1a,8'h1a,8'h1a,8'h3,8'h6,8'h2a,8'h1a,8'h21,8'h6,8'h2a,8'h1a,8'h1a,8'h16,8'h6,8'h6,8'h1b,8'h1a,8'h6,8'h6,8'h6,8'h6,8'h6,8'h6,8'h6,8'h6,8'h9,8'h1a,8'h1a,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h1a,8'h1a,8'h1a,8'h1a,8'h1a,8'h1a,8'h1a,8'h1a,8'ha,8'h6,8'h22,8'h1a,8'h1a,8'h1a,8'h16,8'h7,8'h6,8'h21,8'h1a,8'h1a,8'h2b,8'h2b,8'h1a,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h1a,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h1a,8'h1a,8'h1a,8'h21,8'h6,8'h6,8'h1b,8'h1a,8'h1a,8'h1a,8'h1b,8'h6,8'h6,8'h1b,8'h1a,8'h1a,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h1a,8'h1a,8'h1a,8'h1a,8'h1a,8'h1a,8'h1a,8'h21,8'h6,8'h6,8'h1b,8'h21,8'h6,8'h2a,8'h2b,8'h1a,8'h1a,8'h2b,8'h22,8'h6,8'h21,8'h1a,8'h1a,8'h1a,8'h4,8'h6,8'h2a,8'h1a,8'h21,8'h6,8'h2a,8'h1a,8'h1a,8'h1b,8'h6,8'h6,8'h1b,8'h1a,8'h22,8'h6,8'h3,8'h1a,8'h1a,8'h1a,8'h1a,8'h1a,8'h1a,8'h1a,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h1a,8'h1a,8'h1a,8'h1a,8'h2b,8'h1a,8'h1a,8'h1a,8'h21,8'h6,8'h2a,8'h1a,8'h1a,8'h1a,8'h16,8'h7,8'h6,8'h1b,8'h1a,8'h1a,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h1a,8'h1a,8'h21,8'h6,8'h6,8'h1a,8'h1a,8'h1a,8'h1a,8'h1b,8'h6,8'h6,8'h1b,8'h2b,8'h1a,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h1a,8'h1a,8'h1a,8'h1a,8'h1a,8'h21,8'h6,8'h6,8'h16,8'h21,8'h6,8'h2a,8'h1a,8'h1a,8'h1a,8'h1a,8'h22,8'h6,8'h2,8'h1a,8'h1a,8'h1a,8'h6,8'h6,8'h21,8'h1a,8'h21,8'h6,8'h22,8'h1a,8'h1a,8'h1a,8'h6,8'h6,8'h1b,8'h1a,8'h4,8'h6,8'h9,8'h1a,8'h1a,8'h1a,8'h1a,8'h1a,8'h1a,8'h1a,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h1a,8'h1a,8'h1a,8'h1a,8'h2b,8'h1a,8'h1a,8'h1a,8'h16,8'h6,8'h6,8'h1b,8'h2b,8'h1a,8'h1b,8'h6,8'h6,8'h1a,8'h1a,8'h1a,8'h2b,8'h1a,8'h1a,8'h1a,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h1a,8'h1a,8'h1a,8'h21,8'h6,8'h6,8'h1a,8'h1a,8'h2b,8'h1a,8'h1b,8'h6,8'h6,8'h1b,8'h1a,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h16,8'h6,8'h1b,8'h1a,8'h1a,8'h1a,8'h22,8'h6,8'h3,8'h1a,8'h1b,8'h6,8'h6,8'h1b,8'h2b,8'h2b,8'h2b,8'h1b,8'h6,8'h6,8'h21,8'h1a,8'h3,8'h6,8'h6,8'h1a,8'h1a,8'h21,8'h6,8'h9,8'h1a,8'h1a,8'h1b,8'h6,8'h6,8'h1b,8'h1a,8'h16,8'h6,8'h6,8'h9,8'h1a,8'h1a,8'h2b,8'h2b,8'h1a,8'h1a,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h1a,8'h2b,8'h1a,8'h1a,8'h1a,8'h1a,8'h1a,8'h1a,8'h1a,8'h9,8'h6,8'h2a,8'h1a,8'h16,8'h22,8'h6,8'h21,8'h1a,8'h1a,8'h1a,8'h2b,8'h1a,8'h1a,8'h1a,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h1a,8'h1a,8'h21,8'h6,8'h6,8'h1a,8'h1a,8'h1a,8'h1a,8'h1b,8'h6,8'h6,8'h1b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h16,8'h6,8'h6,8'h6,8'h6,8'h22,8'h6,8'h21,8'h1a,8'h1a,8'h1a,8'h3,8'h6,8'h6,8'h6,8'h6,8'h3,8'h1a,8'h16,8'h6,8'h6,8'h6,8'h6,8'h9,8'h2b,8'h1a,8'h1a,8'h21,8'h6,8'h22,8'h1a,8'h1a,8'h1a,8'h22,8'h6,8'h1b,8'h1a,8'h1a,8'h1a,8'h6,8'h6,8'h6,8'h6,8'h6,8'h6,8'h1a,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h1a,8'h1a,8'h2b,8'h2b,8'h1a,8'h1a,8'h2,8'h6,8'h6,8'h6,8'h6,8'h3,8'h1a,8'h1a,8'h1a,8'h1a,8'h1a,8'h1a,8'h1a,8'h1a,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h1a,8'h1a,8'h1a,8'h21,8'h6,8'h6,8'h1b,8'h1a,8'h2b,8'h1a,8'h1b,8'h6,8'h6,8'h1b,8'h1a,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h1a,8'h1a,8'h1a,8'h1a,8'h1a,8'h1a,8'h1a,8'h1a,8'h1a,8'h1a,8'h1a,8'h1a,8'h1a,8'h1a,8'h1a,8'h2b,8'h2b,8'h1a,8'h1a,8'h1a,8'h1a,8'h1a,8'h1a,8'h1a,8'h1a,8'h1a,8'h1a,8'h1a,8'h1a,8'h1a,8'h1a,8'h1a,8'h1a,8'h2b,8'h1a,8'h1a,8'h2b,8'h1a,8'h1a,8'h1a,8'h2b,8'h1a,8'h2b,8'h2b,8'h1a,8'h2b,8'h1a,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h1a,8'h1a,8'h1a,8'h1a,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h1a,8'h1a,8'h1a,8'h1a,8'h1a,8'h1a,8'h2b,8'h1a,8'h1a,8'h1a,8'h1a,8'h1a,8'h2b,8'h1a,8'h1a,8'h1a,8'h1a,8'h1a,8'h1a,8'h1a,8'h1a,8'h1a,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h1a,8'h1a,8'h1a,8'h2b,8'h1a,8'h1a,8'h1a,8'h1a,8'h1a,8'h1a,8'h1a,8'h1a,8'h1a,8'h2b,8'h2b,8'h1a,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h1a,8'h1a,8'h1a,8'h1a,8'h1a,8'h1a,8'h1a,8'h1a,8'h1a,8'h1a,8'h1a,8'h1a,8'h2b,8'h2b,8'h1a,8'h2b,8'h1a,8'h1a,8'h1a,8'h1a,8'h1a,8'h1a,8'h1a,8'h2b,8'h1a,8'h1a,8'h2b,8'h1a,8'h1a,8'h1a,8'h1a,8'h1a,8'h1a,8'h1a,8'h1a,8'h1a,8'h1a,8'h1a,8'h2b,8'h2b,8'h1a,8'h1a,8'h2b,8'h2b,8'h1a,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h1a,8'h1a,8'h1a,8'h1a,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h1a,8'h1a,8'h1a,8'h1a,8'h1a,8'h1a,8'h2b,8'h1a,8'h1a,8'h1a,8'h1a,8'h2b,8'h1a,8'h1a,8'h1a,8'h2b,8'h1a,8'h1a,8'h1a,8'h1a,8'h1a,8'h1a,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h1a,8'h1a,8'h2b,8'h2b,8'h1a,8'h1a,8'h2b,8'h2b,8'h1a,8'h2b,8'h1a,8'h2b,8'h1a,8'h2b,8'h2b,8'h1a,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h1a,8'h1a,8'h1a,8'h1a,8'h1a,8'h1a,8'h1a,8'h1a,8'h1a,8'h1a,8'h1a,8'h1a,8'h1a,8'h1a,8'h2b,8'h1a,8'h1a,8'h1a,8'h1a,8'h1a,8'h2b,8'h2b,8'h1a,8'h1a,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h1a,8'h1a,8'h1a,8'h1a,8'h1a,8'h1a,8'h1a,8'h1a,8'h1a,8'h2b,8'h2b,8'h2b,8'h2b,8'h1a,8'h2b,8'h2b,8'h2b,8'h2b,8'h1a,8'h1a,8'h1a,8'h1a,8'h2b,8'h2b,8'h1a,8'h1a,8'h1a,8'h2b,8'h2b,8'h1a,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h1a,8'h1a,8'h1a,8'h1a,8'h1a,8'h1a,8'h1a,8'h1a,8'h1a,8'h1a,8'h1a,8'h1a,8'h1a,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h1a,8'h2b,8'h2b,8'h2b,8'h1a,8'h1a,8'h1a,8'h1a,8'h1a,8'h1a,8'h1a,8'h1a,8'h1a,8'h1a,8'h1a,8'h1a,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h1a,8'h1a,8'h1a,8'h1a,8'h1a,8'h1a,8'h1a,8'h1a,8'h1a,8'h2b,8'h1a,8'h1a,8'h1a,8'h1a,8'h2b,8'h2b,8'h1a,8'h1a,8'h2b,8'h2b,8'h1a,8'h1a,8'h1a,8'h1a,8'h2b,8'h2b,8'h1a,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h1a,8'h1a,8'h1a,8'h1a,8'h1a,8'h1a,8'h1a,8'h1a,8'h2b,8'h1a,8'h2b,8'h2b,8'h2b,8'h1a,8'h2b,8'h2b,8'h2b,8'h2b,8'h1a,8'h1a,8'h1a,8'h1a,8'h2b,8'h2b,8'h1a,8'h1a,8'h2b,8'h2b,8'h2b,8'h1a,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h1a,8'h1a,8'h1a,8'h1a,8'h1a,8'h1a,8'h1a,8'h1a,8'h1a,8'h1a,8'h1a,8'h1a,8'h1a,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h1a,8'h2b,8'h2b,8'h2b,8'h1a,8'h1a,8'h1a,8'h1a,8'h1a,8'h1a,8'h1a,8'h1a,8'h1a,8'h1a,8'h1a,8'h1a,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h1a,8'h1a,8'h1a,8'h1a,8'h1a,8'h1a,8'h1a,8'h1a,8'h1a,8'h1a,8'h1a,8'h1a,8'h1a,8'h1a,8'h1a,8'h1a,8'h1a,8'h1a,8'h1a,8'h1a,8'h1a,8'h1a,8'h1a,8'h2b,8'h2b,8'h2b,8'h1a,8'h1a,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h1a,8'h1a,8'h1a,8'h1a,8'h1a,8'h1a,8'h1a,8'h1a,8'h1a,8'h1a,8'h2b,8'h2b,8'h2b,8'h1a,8'h2b,8'h2b,8'h2b,8'h2b,8'h1a,8'h1a,8'h1a,8'h1a,8'h2b,8'h2b,8'h1a,8'h1a,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h1a,8'h1a,8'h1a,8'h1a,8'h1a,8'h1a,8'h1a,8'h2b,8'h1a,8'h1a,8'h1a,8'h1a,8'h1a,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h1a,8'h2b,8'h2b,8'h2b,8'h1a,8'h1a,8'h1a,8'h1a,8'h16,8'h1a,8'h1a,8'h1a,8'h1a,8'h1a,8'h1a,8'h1a,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h1a,8'h1a,8'h1a,8'h1a,8'h1a,8'h1a,8'h1a,8'h1a,8'h1a,8'h2b,8'h1a,8'h1a,8'h1a,8'h1a,8'h2b,8'h2b,8'h1a,8'h1a,8'h2b,8'h1a,8'h1a,8'h1a,8'h1a,8'h2b,8'h2b,8'h2b,8'h1a,8'h1a,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h1a,8'h2b,8'h1a,8'h1a,8'h1a,8'h2b,8'h1a,8'h1a,8'h1a,8'h1a,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h1a,8'h1a,8'h1a,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h1a,8'h1a,8'h1a,8'h1a,8'h1a,8'h1a,8'h1a,8'h1a,8'h1a,8'h1a,8'h1a,8'h1a,8'h1a,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h1a,8'h2b,8'h2b,8'h1a,8'h2b,8'h1a,8'h1a,8'h1a,8'h1a,8'h1a,8'h1a,8'h1a,8'h1a,8'h1a,8'h1a,8'h1a,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h1a,8'h1a,8'h1a,8'h1a,8'h1a,8'h1a,8'h1a,8'h1a,8'h1a,8'h1a,8'h1a,8'h1a,8'h1a,8'h1a,8'h1a,8'h2b,8'h1a,8'h1a,8'h1a,8'h2b,8'h1a,8'h1a,8'h2b,8'h1a,8'h2b,8'h2b,8'h1a,8'h1a,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h1a,8'h1a,8'h2b,8'h2b,8'h1a,8'h1a,8'h1a,8'h1a,8'h2b,8'h1a,8'h2b,8'h2b,8'h2b,8'h1a,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h1a,8'h1a,8'h1a,8'h1a,8'h1a,8'h1a,8'h2b,8'h1a,8'h1a,8'h1a,8'h1a,8'h1a,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h1a,8'h2b,8'h2b,8'h2b,8'h2b,8'h1a,8'h1a,8'h1a,8'h1a,8'h1a,8'h1a,8'h1a,8'h1a,8'h1a,8'h1a,8'h1a,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h1a,8'h1a,8'h1a,8'h1a,8'h1a,8'h1a,8'h1a,8'h1a,8'h2b,8'h2b,8'h1a,8'h1a,8'h1a,8'h1a,8'h1a,8'h2b,8'h1a,8'h1a,8'h1a,8'h1a,8'h1a,8'h1a,8'h2b,8'h2b,8'h2b,8'h1a,8'h1a,8'h1a,8'h2b,8'h2b,8'h2b,8'h1a,8'h2b,8'h2b,8'h1a,8'h2b,8'h2b,8'h2b,8'h1a,8'h1a,8'h1a,8'h2b,8'h1a,8'h1a,8'h2b,8'h2b,8'h2b,8'h1a,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h1a,8'h1a,8'h1a,8'h1a,8'h1a,8'h1a,8'h1a,8'h1a,8'h1a,8'h1a,8'h1a,8'h1a,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h1a,8'h2b,8'h2b,8'h2b,8'h2b,8'h1a,8'h1a,8'h1a,8'h1a,8'h1a,8'h1a,8'h1a,8'h1a,8'h1a,8'h1a,8'h1a,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h1a,8'h1a,8'h1a,8'h1a,8'h1a,8'h1a,8'h1a,8'h1a,8'h1a,8'h1a,8'h21,8'h6,8'h6,8'h6,8'h6,8'h6,8'h6,8'h1b,8'h1a,8'h1a,8'h1a,8'h1a,8'h1a,8'h1a,8'h1a,8'h1a,8'h1a,8'h1a,8'h2b,8'h2b,8'h2b,8'h1a,8'h1a,8'h1a,8'h1a,8'h1a,8'h2b,8'h2b,8'h1a,8'h1a,8'h1a,8'h2b,8'h1a,8'h1a,8'h2b,8'h2b,8'h1a,8'h1a,8'h1a,8'h1a,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h1a,8'h1a,8'h1a,8'h2b,8'h1a,8'h1a,8'h1a,8'h1a,8'h9,8'h6,8'h2a,8'h1a,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h1a,8'h2b,8'h2b,8'h2b,8'h2b,8'h1a,8'h1a,8'h1a,8'h16,8'h6,8'h6,8'h1a,8'h1a,8'h1a,8'h1a,8'h1a,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h1a,8'h1a,8'h1a,8'h1a,8'h1a,8'h1a,8'h1a,8'h1a,8'h1a,8'h2b,8'h21,8'h6,8'h9,8'h1a,8'h1a,8'h21,8'h6,8'h6,8'h21,8'h1a,8'h1a,8'h1a,8'h1a,8'h1a,8'h1a,8'h1a,8'h1a,8'h1a,8'h2b,8'h2b,8'h2b,8'h1a,8'h1a,8'h1a,8'h1a,8'h1a,8'h2b,8'h1a,8'h1a,8'h1a,8'h2b,8'h2b,8'h1a,8'h1a,8'h2b,8'h2b,8'h1a,8'h1a,8'h1a,8'h1a,8'h2b,8'h2b,8'h2b,8'h1a,8'h1a,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h1a,8'h2b,8'h2b,8'h2b,8'h1a,8'h1a,8'h1a,8'h2b,8'h1a,8'h1a,8'h1a,8'h1a,8'h9,8'h6,8'h2a,8'h1a,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h1a,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h1a,8'h1a,8'h1b,8'h6,8'h6,8'h1a,8'h1a,8'h1a,8'h1a,8'h1a,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h1a,8'h1a,8'h1a,8'h1a,8'h2b,8'h1a,8'h1a,8'h1a,8'h2b,8'h2b,8'h21,8'h6,8'h6,8'h1a,8'h1a,8'h2b,8'h3,8'h6,8'h6,8'h1a,8'h1a,8'h1a,8'h1a,8'h1a,8'h1a,8'h1a,8'h1a,8'h1a,8'h2b,8'h1a,8'h2b,8'h1a,8'h1a,8'h1a,8'h1a,8'h1a,8'h1a,8'h1a,8'h1a,8'h1a,8'h2b,8'h1a,8'h1a,8'h1a,8'h1a,8'h2b,8'h1a,8'h1a,8'h1a,8'h1a,8'h1a,8'h2b,8'h1a,8'h1a,8'h1a,8'h1a,8'h2b,8'h2b,8'h1a,8'h1a,8'h2b,8'h2b,8'h2b,8'h1a,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h1a,8'h2b,8'h2b,8'h2b,8'h1a,8'h1a,8'h1a,8'h2b,8'h1a,8'h1a,8'h1a,8'h1a,8'h9,8'h6,8'h2a,8'h1a,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h1a,8'h2b,8'h1a,8'h2b,8'h2b,8'h1a,8'h1a,8'h1a,8'h1b,8'h6,8'h6,8'h1a,8'h1a,8'h1a,8'h1a,8'h1a,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h1a,8'h1a,8'h1a,8'h1a,8'h2b,8'h1a,8'h1a,8'h1a,8'h1a,8'h1a,8'h21,8'h6,8'h9,8'h1a,8'h1a,8'h1a,8'h21,8'h6,8'h6,8'h1a,8'h1b,8'h6,8'h6,8'h6,8'h6,8'h6,8'h1b,8'h1a,8'h1a,8'h21,8'h6,8'h6,8'h6,8'h6,8'h6,8'h22,8'h1a,8'h1a,8'h1a,8'h1a,8'h1a,8'h6,8'h6,8'h6,8'h6,8'h6,8'h1b,8'h1a,8'h1a,8'h21,8'h6,8'h6,8'h6,8'h6,8'h6,8'h3,8'h2b,8'h2b,8'h1a,8'h1a,8'h1a,8'h2b,8'h2b,8'h1a,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h1a,8'h2b,8'h2b,8'h2b,8'h1a,8'h1a,8'h1a,8'h2b,8'h1a,8'h1a,8'h1a,8'h1a,8'h9,8'h6,8'h2a,8'h1a,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h1a,8'h1a,8'h1a,8'h2b,8'h1a,8'h1a,8'h21,8'h6,8'h6,8'h1a,8'h2b,8'h1a,8'h1a,8'h1a,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h1a,8'h1a,8'h1a,8'h1a,8'h1a,8'h1a,8'h1a,8'h2b,8'h2b,8'h1a,8'h1,8'h6,8'h22,8'h1a,8'h2b,8'h2b,8'h3,8'h6,8'h6,8'h1a,8'h1a,8'h1a,8'h1a,8'h1a,8'ha,8'h6,8'h22,8'h1b,8'h2b,8'h21,8'h6,8'h9,8'h1a,8'h1a,8'h9,8'h6,8'h6,8'h1a,8'h1a,8'h1a,8'h6,8'h6,8'h21,8'h1a,8'h21,8'h6,8'h6,8'h1b,8'h1a,8'h21,8'h6,8'h22,8'h1a,8'h1a,8'h1a,8'h1a,8'h2b,8'h1a,8'h1a,8'h1a,8'h1a,8'h2b,8'h1a,8'h1a,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h1a,8'h1a,8'h2b,8'h2b,8'h2b,8'h1a,8'h2b,8'h2b,8'h1a,8'h1a,8'h1a,8'h1a,8'h9,8'h6,8'h2a,8'h1a,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h1a,8'h1a,8'h1a,8'h1a,8'h2b,8'h1a,8'h1a,8'h16,8'h6,8'h6,8'h1a,8'h1a,8'h1a,8'h1a,8'h1a,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h1a,8'h1a,8'h1a,8'h1a,8'h1a,8'h1a,8'h1a,8'h2b,8'h2b,8'h1a,8'h21,8'h6,8'h9,8'h1a,8'h1a,8'h21,8'h6,8'h6,8'h21,8'h2b,8'h1a,8'h1a,8'h1a,8'h1a,8'h16,8'h6,8'h6,8'h1b,8'h1a,8'h21,8'h6,8'h22,8'h1a,8'h1a,8'h18,8'h6,8'h6,8'h3,8'h1a,8'ha,8'h6,8'h2a,8'h1a,8'h1a,8'h1a,8'h3,8'h6,8'h21,8'h1a,8'h21,8'h6,8'h6,8'h1a,8'h1a,8'h1a,8'h1a,8'h2b,8'h1a,8'h1a,8'h1a,8'h1a,8'h2b,8'h1a,8'h1a,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h1a,8'h1a,8'h2b,8'h2b,8'h2b,8'h1a,8'h2b,8'h2b,8'h1a,8'h1a,8'h1a,8'h1a,8'h9,8'h6,8'h2a,8'h1a,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h1a,8'h1a,8'h1a,8'h1a,8'h2b,8'h2b,8'h1a,8'h1a,8'h1b,8'h6,8'h6,8'h1a,8'h1a,8'h1a,8'h1a,8'h1a,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h1a,8'h1a,8'h1a,8'h1a,8'h1a,8'h1a,8'h1a,8'h2b,8'h2b,8'h1a,8'h0,8'h6,8'h6,8'h6,8'h6,8'h6,8'h6,8'h16,8'h1a,8'h1a,8'h1a,8'h9,8'h6,8'h6,8'h6,8'h6,8'h6,8'h1a,8'h1a,8'h4,8'h6,8'h2a,8'h1a,8'h1a,8'h18,8'h9,8'h6,8'h2a,8'h1a,8'h6,8'h6,8'h6,8'h6,8'h6,8'h6,8'h6,8'h6,8'h2,8'h1a,8'h21,8'h6,8'h22,8'h1a,8'h1a,8'h1a,8'h1a,8'h2b,8'h1a,8'h1a,8'h1a,8'h1a,8'h2b,8'h1a,8'h1a,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h1a,8'h1a,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h1a,8'h1a,8'h1a,8'h1a,8'h9,8'h6,8'h2a,8'h1a,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h1a,8'h2b,8'h1a,8'h1a,8'h1a,8'h1a,8'h1a,8'h1a,8'h1b,8'h6,8'h6,8'h1a,8'h1a,8'h1a,8'h1a,8'h1a,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h1a,8'h1a,8'h1a,8'h1a,8'h1a,8'h1a,8'h1a,8'h2b,8'h1a,8'h1a,8'h0,8'h6,8'h9,8'h1a,8'h1a,8'h1a,8'h2b,8'h1a,8'h1a,8'h1a,8'h6,8'h6,8'h2a,8'h1a,8'h16,8'h6,8'h6,8'h1b,8'h1a,8'h1b,8'h6,8'h2a,8'h1a,8'h1a,8'h1a,8'h9,8'h6,8'h2a,8'h1a,8'h6,8'h6,8'h3,8'h1a,8'h1a,8'h1a,8'h2b,8'h1a,8'h1a,8'h1a,8'h21,8'h6,8'h6,8'h1a,8'h1a,8'h1a,8'h1a,8'h2b,8'h1a,8'h1a,8'h1a,8'h1a,8'h2b,8'h1a,8'h1a,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h1a,8'h1a,8'h2b,8'h2b,8'h2b,8'h1a,8'h2b,8'h2b,8'h1a,8'h1a,8'h1a,8'h1a,8'h9,8'h6,8'h2a,8'h1a,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h1a,8'h1a,8'h1a,8'h2b,8'h2b,8'h1a,8'h1a,8'h16,8'h6,8'h6,8'h1a,8'h2b,8'h1a,8'h1a,8'h1a,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h1a,8'h1a,8'h1a,8'h1a,8'h1a,8'h1a,8'h1a,8'h2b,8'h1a,8'h1a,8'h21,8'h6,8'h22,8'h1a,8'h1a,8'h1a,8'h2b,8'h1a,8'h1a,8'h1b,8'h6,8'h6,8'h1a,8'h1a,8'h16,8'h22,8'h6,8'h1b,8'h1a,8'h21,8'h6,8'h2a,8'h1a,8'h1a,8'h18,8'h22,8'h6,8'h21,8'h1a,8'ha,8'h6,8'h2a,8'h1a,8'h1a,8'h1a,8'h2b,8'h1a,8'h1a,8'h18,8'h21,8'h6,8'h22,8'h1a,8'h1a,8'h1a,8'h1a,8'h2b,8'h1a,8'h1a,8'h1a,8'h1a,8'h2b,8'h1a,8'h1a,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h1a,8'h1a,8'h1a,8'h2b,8'h2b,8'h1a,8'h2b,8'h2b,8'h1a,8'h1a,8'h1a,8'h1a,8'h9,8'h6,8'h2a,8'h1a,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h1a,8'h1a,8'h1a,8'h1a,8'h1a,8'h1a,8'h1a,8'h1a,8'h21,8'h6,8'h2a,8'h1a,8'h1a,8'h1a,8'h1a,8'h1a,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h1a,8'h1a,8'h1a,8'h1a,8'h1a,8'h1a,8'h1a,8'h2b,8'h2b,8'h1a,8'h21,8'h6,8'h22,8'h1a,8'h1a,8'h1a,8'h1a,8'h1a,8'h1a,8'h1a,8'h6,8'h6,8'h3,8'h1a,8'h16,8'h6,8'h6,8'h1b,8'h1a,8'h21,8'h6,8'h6,8'h1a,8'h1a,8'ha,8'h6,8'h6,8'h1a,8'h18,8'h18,8'h6,8'h6,8'h2a,8'h1a,8'h1a,8'h1a,8'h1a,8'h1a,8'h1a,8'h21,8'h6,8'h6,8'h1a,8'h1a,8'h1a,8'h1a,8'h2b,8'h1a,8'h1a,8'h1a,8'h1a,8'h2b,8'h1a,8'h1a,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h1a,8'h1a,8'h1a,8'h2b,8'h2b,8'h1a,8'h1a,8'h2b,8'h1a,8'h1a,8'h1a,8'h1a,8'h9,8'h6,8'h2a,8'h1a,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h1a,8'h1a,8'h1a,8'h3,8'h6,8'h21,8'h1a,8'h16,8'h6,8'h6,8'h21,8'h1a,8'h2b,8'h1a,8'h1a,8'h1a,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h1a,8'h1a,8'h2b,8'h1a,8'h21,8'h6,8'h22,8'h1a,8'h1a,8'h1a,8'h1a,8'h1a,8'h1a,8'h1a,8'h1b,8'h22,8'h6,8'h6,8'h6,8'h6,8'h6,8'h1b,8'h1a,8'h21,8'h6,8'h6,8'h6,8'h6,8'h6,8'h22,8'h16,8'h1a,8'h2b,8'h1a,8'h1a,8'h22,8'h6,8'h6,8'h6,8'h6,8'h6,8'h1a,8'h1a,8'h21,8'h6,8'h6,8'h1b,8'h1a,8'h1a,8'h1a,8'h1a,8'h2b,8'h1a,8'h1a,8'h1a,8'h1a,8'h2b,8'h1a,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h1a,8'h2b,8'h1a,8'h3,8'h6,8'h9,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h1a,8'h1a,8'h1a,8'h1a,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h1a,8'h1a,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h1a,8'h2b,8'h2b,8'h1a,8'h3,8'h6,8'h6,8'h6,8'h22,8'h1b,8'h1a,8'h1a,8'h1a,8'h2b,8'h1a,8'h1a,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h1a,8'h1a,8'h2b,8'h1a,8'h1a,8'h1a,8'h1a,8'h1a,8'h1a,8'h1a,8'h1a,8'h1a,8'h1a,8'h1a,8'h1a,8'h1a,8'h2b,8'h2b,8'h1a,8'h2b,8'h1a,8'h1a,8'h1a,8'h21,8'h6,8'h2a,8'h1a,8'h1a,8'h1a,8'h1a,8'h1a,8'h1a,8'h1a,8'h1a,8'h1a,8'h1a,8'h1a,8'h1a,8'h1a,8'h1a,8'h1a,8'h1a,8'h1a,8'h2b,8'h1a,8'h1a,8'h1a,8'h1a,8'h1a,8'h1a,8'h1a,8'h2b,8'h1a,8'h1a,8'h1a,8'h1a,8'h2b,8'h1a,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h1a,8'h2b,8'h1a,8'h1a,8'h1a,8'h1a,8'h1a,8'h1a,8'h2b,8'h2b,8'h2b,8'h2b,8'h1a,8'h1a,8'h1a,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h1a,8'h1a,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h1a,8'h1a,8'h1a,8'h1a,8'h1a,8'h1a,8'h1a,8'h2b,8'h1a,8'h2b,8'h1a,8'h1a,8'h2b,8'h2b,8'h1a,8'h1a,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h1a,8'h1a,8'h1a,8'h1a,8'h2b,8'h2b,8'h2b,8'h1a,8'h1a,8'h1a,8'h1a,8'h1a,8'h1a,8'h1a,8'h1a,8'h1a,8'h2b,8'h1a,8'h1a,8'h1a,8'h2b,8'h1a,8'h1a,8'h21,8'h6,8'h2a,8'h1a,8'h1a,8'h1a,8'h1a,8'h1a,8'h1a,8'h1a,8'h2b,8'h1a,8'h2b,8'h1a,8'h1a,8'h1a,8'h1a,8'h1a,8'h1a,8'h1a,8'h2b,8'h1a,8'h1a,8'h1a,8'h1a,8'h2b,8'h2b,8'h2b,8'h2b,8'h1a,8'h1a,8'h1a,8'h1a,8'h2b,8'h1a,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h1a,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h1a,8'h2b,8'h2b,8'h2b,8'h2b,8'h1a,8'h1a,8'h1a,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h1a,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h1a,8'h2b,8'h1a,8'h1a,8'h1a,8'h1a,8'h1a,8'h1a,8'h2b,8'h2b,8'h1a,8'h1a,8'h2b,8'h1a,8'h1a,8'h1a,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h1a,8'h1a,8'h1a,8'h2b,8'h1a,8'h1a,8'h1a,8'h2b,8'h1a,8'h1a,8'h1a,8'h1a,8'h1a,8'h1a,8'h1a,8'h2b,8'h2b,8'h2b,8'h2b,8'h1a,8'h2b,8'h1a,8'h1a,8'h21,8'h6,8'h2a,8'h1a,8'h2b,8'h1a,8'h1a,8'h1a,8'h1a,8'h1a,8'h1a,8'h2b,8'h2b,8'h1a,8'h1a,8'h1a,8'h1a,8'h1a,8'h1a,8'h1a,8'h1a,8'h1a,8'h2b,8'h1a,8'h1a,8'h2b,8'h1a,8'h2b,8'h2b,8'h1a,8'h1a,8'h1a,8'h1a,8'h2b,8'h1a,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h1a,8'h1a,8'h1a,8'h1a,8'h1a,8'h1a,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h1a,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h1a,8'h2b,8'h2b,8'h1a,8'h1a,8'h1a,8'h1a,8'h2b,8'h1a,8'h1a,8'h1a,8'h2b,8'h1a,8'h1a,8'h1a,8'h1a,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h1a,8'h1a,8'h1a,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h1a,8'h1a,8'h1a,8'h1a,8'h1a,8'h1a,8'h1a,8'h1a,8'h1a,8'h2b,8'h1a,8'h1a,8'h2b,8'h1a,8'h1a,8'h1a,8'h1a,8'h1a,8'h1a,8'h1a,8'h1a,8'h1a,8'h1a,8'h1a,8'h2b,8'h2b,8'h1a,8'h2b,8'h1a,8'h1a,8'h1a,8'h1a,8'h1a,8'h1a,8'h1a,8'h2b,8'h1a,8'h2b,8'h1a,8'h1a,8'h2b,8'h2b,8'h2b,8'h2b,8'h1a,8'h1a,8'h2b,8'h1a,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h1a,8'h2b,8'h2b,8'h1a,8'h1a,8'h2b,8'h2b,8'h1a,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h1a,8'h2b,8'h1a,8'h1a,8'h1a,8'h1a,8'h1a,8'h1a,8'h2b,8'h2b,8'h1a,8'h1a,8'h1a,8'h2b,8'h2b,8'h1a,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h1a,8'h1a,8'h1a,8'h1a,8'h1a,8'h2b,8'h2b,8'h1a,8'h1a,8'h2b,8'h2b,8'h1a,8'h1a,8'h1a,8'h1a,8'h1a,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h1a,8'h1a,8'h1a,8'h1a,8'h1a,8'h2b,8'h2b,8'h2b,8'h1a,8'h1a,8'h1a,8'h2b,8'h2b,8'h2b,8'h1a,8'h1a,8'h1a,8'h1a,8'h1a,8'h1a,8'h1a,8'h2b,8'h2b,8'h1a,8'h1a,8'h2b,8'h1a,8'h2b,8'h2b,8'h2b,8'h2b,8'h1a,8'h2b,8'h1a,8'h1a,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h1a,8'h2b,8'h2b,8'h2b,8'h1a,8'h1a,8'h1a,8'h1a,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h1a,8'h1a,8'h1a,8'h1a,8'h1a,8'h1a,8'h1a,8'h1a,8'h2b,8'h1a,8'h1a,8'h1a,8'h1a,8'h2b,8'h1a,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h1a,8'h1a,8'h1a,8'h1a,8'h1a,8'h1a,8'h2b,8'h1a,8'h1a,8'h2b,8'h1a,8'h1a,8'h1a,8'h1a,8'h1a,8'h1a,8'h2b,8'h1a,8'h1a,8'h2b,8'h1a,8'h1a,8'h1a,8'h1a,8'h1a,8'h1a,8'h1a,8'h2b,8'h2b,8'h1a,8'h1a,8'h1a,8'h1a,8'h1a,8'h1a,8'h2b,8'h1a,8'h1a,8'h1a,8'h1a,8'h1a,8'h1a,8'h1a,8'h1a,8'h2b,8'h1a,8'h1a,8'h2b,8'h1a,8'h1a,8'h1a,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h1a,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h1a,8'h1a,8'h1a,8'h2b,8'h2b,8'h2b,8'h2b,8'h1a,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h1a,8'h1a,8'h1a,8'h1a,8'h1a,8'h1a,8'h1a,8'h1a,8'h2b,8'h1a,8'h1a,8'h1a,8'h2b,8'h2b,8'h1a,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h1a,8'h1a,8'h1a,8'h1a,8'h1a,8'h1a,8'h1a,8'h2b,8'h1a,8'h2b,8'h2b,8'h1a,8'h1a,8'h1a,8'h1a,8'h1a,8'h1a,8'h1a,8'h2b,8'h1a,8'h2b,8'h2b,8'h1a,8'h1a,8'h1a,8'h1a,8'h1a,8'h1a,8'h2b,8'h1a,8'h2b,8'h1a,8'h2b,8'h1a,8'h2b,8'h1a,8'h2b,8'h1a,8'h1a,8'h1a,8'h2b,8'h1a,8'h1a,8'h2b,8'h1a,8'h1a,8'h1a,8'h1a,8'h1a,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h1a,8'h1a,8'h1a,8'h1a,8'h2b,8'h2b,8'h1a,8'h1a,8'h2b,8'h2b,8'h1a,8'h1a,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h1a,8'h1a,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h1a,8'h2b,8'h2b,8'h1a,8'h1a,8'h1a,8'h1a,8'h1a,8'h2b,8'h2b,8'h1a,8'h1a,8'h1a,8'h2b,8'h1a,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h1a,8'h1a,8'h1a,8'h1a,8'h1a,8'h1a,8'h1a,8'h1a,8'h2b,8'h2b,8'h1a,8'h1a,8'h1a,8'h1a,8'h1a,8'h1a,8'h1a,8'h2b,8'h1a,8'h2b,8'h2b,8'h1a,8'h1a,8'h1a,8'h1a,8'h1a,8'h1a,8'h1a,8'h1a,8'h2b,8'h2b,8'h1a,8'h2b,8'h1a,8'h1a,8'h2b,8'h1a,8'h1a,8'h2b,8'h2b,8'h2b,8'h1a,8'h1a,8'h2b,8'h1a,8'h1a,8'h1a,8'h2b,8'h2b,8'h1a,8'h2b,8'h2b,8'h2b,8'h1a,8'h2b,8'h1a,8'h1a,8'h2b,8'h1a,8'h1a,8'h1a,8'h1a,8'h1a,8'h2b,8'h1a,8'h1a,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h1a,8'h1a,8'h1a,8'h1a,8'h2b,8'h2b,8'h2b,8'h1a,8'h2b,8'h1a,8'h1a,8'h1a,8'h2b,8'h1a,8'h2b,8'h1a,8'h1a,8'h2b,8'h2b,8'h1a,8'h1a,8'h1a,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h1a,8'h1a,8'h1a,8'h1a,8'h1a,8'h1a,8'h1a,8'h1a,8'h2b,8'h2b,8'h1a,8'h1a,8'h1a,8'h1a,8'h1a,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h1a,8'h1a,8'h1a,8'h1a,8'h1a,8'h1a,8'h1a,8'h3,8'h6,8'h6,8'h6,8'h6,8'h6,8'h1b,8'h1a,8'h1a,8'h1a,8'h2b,8'h1a,8'h2b,8'h1a,8'h2b,8'h1a,8'h1a,8'h9,8'h6,8'h9,8'h1a,8'h1a,8'h1a,8'h2b,8'h2b,8'h2b,8'h1a,8'h1a,8'h1a,8'h1a,8'h1a,8'h2b,8'h1a,8'h1a,8'h1a,8'h1a,8'h1a,8'h1a,8'h1a,8'h2b,8'h2b,8'h1a,8'h1a,8'h2b,8'h1a,8'h1a,8'h2b,8'h2b,8'h2b,8'h1a,8'h1a,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h1a,8'h1a,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h1a,8'h1a,8'h1a,8'h1a,8'h1a,8'h1a,8'h2b,8'h6,8'h6,8'h6,8'h6,8'h6,8'h9,8'h16,8'h2b,8'h1a,8'h1a,8'h1a,8'h1a,8'h2b,8'h1a,8'h1a,8'h1a,8'h1a,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h1a,8'h2b,8'h1a,8'h1a,8'h1a,8'h1a,8'h3,8'h6,8'h22,8'h1a,8'h1a,8'h1a,8'h6,8'h6,8'h6,8'h1a,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h1a,8'h1a,8'h1a,8'h1a,8'h1a,8'h1a,8'h9,8'h6,8'h9,8'h2b,8'h1a,8'h2b,8'h21,8'h1b,8'h1a,8'h1a,8'h2b,8'h1a,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h1a,8'hb,8'h6,8'h2,8'h1a,8'h1a,8'h1a,8'h1a,8'h2b,8'h1a,8'h2b,8'h1a,8'h1a,8'h1a,8'h2b,8'h1a,8'h2b,8'h1a,8'h2b,8'h1a,8'h1a,8'h1a,8'h1a,8'h1a,8'h1a,8'h1a,8'h1a,8'h1a,8'h2b,8'h2b,8'h2b,8'h1a,8'h1a,8'h1a,8'h1a,8'h1a,8'h2b,8'h1a,8'h1a,8'h1a,8'h1a,8'h2b,8'h2b,8'h2b,8'h1a,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h1a,8'h2b,8'h2b,8'h2b,8'h2b,8'h1a,8'h1a,8'h1a,8'h1a,8'h1a,8'h21,8'h6,8'h6,8'h3,8'h1a,8'h1a,8'h9,8'h6,8'h6,8'h16,8'h2b,8'h1a,8'h1a,8'h1a,8'h1a,8'h1a,8'h1a,8'h1a,8'h1a,8'h1a,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h1a,8'h2b,8'h1a,8'h1a,8'h1a,8'h1a,8'h3,8'h6,8'h22,8'h2b,8'h1a,8'h6,8'h6,8'h22,8'h1a,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h1a,8'h1a,8'h1a,8'h1a,8'h1a,8'h1b,8'h6,8'h6,8'h21,8'h1a,8'h2b,8'h1a,8'h1a,8'h1a,8'h1a,8'h1a,8'h1a,8'h2b,8'h1a,8'h2b,8'h2b,8'h2b,8'h1a,8'h1a,8'h1a,8'h1a,8'h1a,8'h1a,8'h1a,8'h1a,8'h1a,8'h2b,8'h1a,8'h1a,8'h1a,8'h1a,8'h1a,8'h1a,8'h1a,8'h2b,8'h2b,8'h1a,8'h1a,8'h1a,8'h1a,8'h1a,8'h1a,8'h1a,8'h1a,8'h1a,8'h2b,8'h1a,8'h1a,8'h1a,8'h1a,8'h1a,8'h1a,8'h1a,8'h1a,8'h2b,8'h2b,8'h2b,8'h2b,8'h1a,8'h1a,8'h1a,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h1a,8'h1a,8'h2b,8'h2b,8'h2b,8'h1a,8'h1a,8'h1a,8'h1a,8'h16,8'h6,8'h6,8'h3,8'h2b,8'h1a,8'h1a,8'h1a,8'h3,8'h6,8'h22,8'h2b,8'h1a,8'h1a,8'h1a,8'h1a,8'h1a,8'h1a,8'h1a,8'h1a,8'h1a,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h1a,8'h2b,8'h2b,8'h1a,8'h1a,8'h1a,8'h4,8'h6,8'h9,8'h1a,8'h9,8'h6,8'h9,8'h1a,8'h1a,8'h1a,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h1a,8'h1a,8'h1a,8'h1a,8'h1a,8'h1a,8'h22,8'h6,8'h9,8'h1a,8'h1a,8'h1a,8'h1a,8'h1a,8'h1a,8'h1a,8'h2b,8'h3,8'h6,8'h6,8'h6,8'h6,8'h6,8'h21,8'h9,8'h6,8'h9,8'h1a,8'h16,8'h6,8'h6,8'h6,8'h6,8'h6,8'h1b,8'h1a,8'h1b,8'h22,8'h6,8'h6,8'h6,8'h6,8'h1b,8'h1a,8'h1a,8'h16,8'h6,8'h6,8'h6,8'h6,8'h22,8'h1a,8'h1a,8'h1a,8'h21,8'h6,8'h6,8'h6,8'h6,8'h6,8'h21,8'h1b,8'h2b,8'h2b,8'h2b,8'h1a,8'h1a,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h1a,8'h1a,8'h2b,8'h2b,8'h2b,8'h1a,8'h1a,8'h1a,8'h1a,8'h3,8'h6,8'h6,8'h1a,8'h1a,8'h1a,8'h1a,8'h1a,8'h1a,8'h22,8'h6,8'h21,8'h1a,8'h1a,8'h1a,8'h1a,8'h1a,8'h1a,8'h1a,8'h1a,8'h1a,8'h2b,8'h1a,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h1a,8'h2b,8'h1a,8'h1a,8'h1a,8'h1a,8'h3,8'h6,8'h22,8'h9,8'h6,8'h6,8'h1a,8'h1a,8'h1a,8'h1a,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h1a,8'h2b,8'h1a,8'h1a,8'h1a,8'h1a,8'h1a,8'h1a,8'h21,8'h6,8'h6,8'h6,8'h6,8'h6,8'h1b,8'h1a,8'h1a,8'h1a,8'h6,8'h6,8'h9,8'h1a,8'h2b,8'h2b,8'h1a,8'h1a,8'h9,8'h6,8'h9,8'h1a,8'h9,8'h6,8'h3,8'h1a,8'h1a,8'h1a,8'h1a,8'h1a,8'h9,8'h6,8'h3,8'h1a,8'h1a,8'h1a,8'h1a,8'h1a,8'h16,8'h6,8'h6,8'h21,8'h1a,8'ha,8'h6,8'h6,8'h1a,8'h2b,8'h21,8'h6,8'h6,8'h1a,8'h1a,8'h1a,8'h1a,8'h2b,8'h2b,8'h1a,8'h1a,8'h1a,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h1a,8'h1a,8'h2b,8'h2b,8'h2b,8'h1a,8'h1a,8'h1a,8'h1a,8'h9,8'h6,8'h9,8'h1a,8'h1a,8'h1a,8'h1a,8'h1a,8'h16,8'h6,8'h6,8'h21,8'h1a,8'h1a,8'h1a,8'h1a,8'h1a,8'h1a,8'h1a,8'h1a,8'h1a,8'h2b,8'h1a,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h1a,8'h2b,8'h1a,8'h1a,8'h1a,8'h1a,8'h4,8'h6,8'h6,8'h6,8'h6,8'h1b,8'h1a,8'h1a,8'h1a,8'h1a,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h1a,8'h2b,8'h1a,8'h2b,8'h1a,8'h1a,8'h1a,8'h1a,8'h1a,8'h1a,8'h1a,8'h1b,8'h22,8'h6,8'h6,8'h6,8'h6,8'h2,8'h1a,8'h21,8'h6,8'h9,8'h1a,8'h2b,8'h1a,8'h2b,8'h2b,8'h1a,8'h9,8'h6,8'h2,8'h1a,8'h6,8'h6,8'h21,8'h1a,8'h1a,8'h2b,8'h1a,8'h1a,8'h6,8'h6,8'h21,8'h1a,8'h2b,8'h2b,8'h1a,8'h1a,8'h9,8'h6,8'h2a,8'h1a,8'h1a,8'h18,8'h22,8'h6,8'h21,8'h1a,8'h21,8'h6,8'h6,8'h1a,8'h1a,8'h1a,8'h2b,8'h2b,8'h1a,8'h1a,8'h2b,8'h2b,8'h2b,8'h1a,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h1a,8'h1a,8'h2b,8'h2b,8'h2b,8'h1a,8'h1a,8'h1a,8'h1a,8'h9,8'h6,8'h9,8'h2b,8'h2b,8'h1a,8'h1a,8'h1a,8'h1a,8'h6,8'h6,8'h2a,8'h1a,8'h1a,8'h1a,8'h1a,8'h1a,8'h1a,8'h1a,8'h1a,8'h1a,8'h1a,8'h1a,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h1a,8'h1a,8'h2b,8'h1a,8'h1a,8'h1a,8'h3,8'h6,8'h6,8'h6,8'h2,8'h1a,8'h1a,8'h1a,8'h1a,8'h1a,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h1a,8'h2b,8'h1a,8'h2b,8'h1a,8'h1a,8'h1a,8'h1a,8'h1a,8'h1a,8'h1a,8'h1a,8'h1a,8'h1a,8'h1a,8'h22,8'h6,8'h6,8'h16,8'h9,8'h6,8'h9,8'h2b,8'h1a,8'h1a,8'h2b,8'h1a,8'h1a,8'h9,8'h6,8'h9,8'h1a,8'h21,8'h6,8'h6,8'h6,8'h1b,8'h1a,8'h1a,8'h1a,8'h21,8'h6,8'h6,8'h6,8'h21,8'h1a,8'h1a,8'h1a,8'h22,8'h6,8'h21,8'h1a,8'h1a,8'h1a,8'h3,8'h6,8'h2,8'h1a,8'h21,8'h6,8'h6,8'h1a,8'h1a,8'h1a,8'h1a,8'h2b,8'h2b,8'h2b,8'h2b,8'h1a,8'h1a,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h1a,8'h1a,8'h2b,8'h2b,8'h2b,8'h1a,8'h1a,8'h1a,8'h1a,8'h9,8'h6,8'h9,8'h1a,8'h1a,8'h1a,8'h1a,8'h1a,8'h1a,8'h6,8'h6,8'h21,8'h1a,8'h1a,8'h1a,8'h1a,8'h1a,8'h1a,8'h1a,8'h1a,8'h1a,8'h1a,8'h1a,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h1a,8'h2b,8'h1a,8'h1a,8'h1a,8'h1a,8'h3,8'h6,8'h6,8'h6,8'h6,8'h22,8'h1a,8'h1a,8'h1a,8'h1a,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h1a,8'h2b,8'h1a,8'h1a,8'h1a,8'h1a,8'h2b,8'h1a,8'h1a,8'h1a,8'h1a,8'h1a,8'h1a,8'h1a,8'h1a,8'h1a,8'h1a,8'h1a,8'h1a,8'h1a,8'h2b,8'h1a,8'h1a,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h1a,8'h1a,8'h1a,8'h1a,8'h1a,8'h1a,8'h1a,8'h1a,8'h1a,8'h21,8'h6,8'h6,8'h1b,8'h9,8'h6,8'h2a,8'h1a,8'h1a,8'h1a,8'h2b,8'h1a,8'h1a,8'h9,8'h6,8'h2,8'h1a,8'h1a,8'h1a,8'h3,8'h6,8'h6,8'h6,8'h16,8'h1a,8'h2b,8'h1a,8'h21,8'h6,8'h6,8'h6,8'h1b,8'h1a,8'h22,8'h6,8'h21,8'h1a,8'h1a,8'h1a,8'h3,8'h6,8'h2a,8'h2b,8'h21,8'h6,8'h6,8'h1a,8'h1a,8'h1a,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h1a,8'h1a,8'h1a,8'h3,8'h6,8'h6,8'h1a,8'h1a,8'h1a,8'h2b,8'h1a,8'h1a,8'h6,8'h6,8'h21,8'h1a,8'h1a,8'h1a,8'h1a,8'h1a,8'h1a,8'h1a,8'h1a,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h1a,8'h1a,8'h1a,8'h1a,8'h2b,8'ha,8'h6,8'h22,8'h1a,8'h6,8'h6,8'h22,8'h1a,8'h1a,8'h1a,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h1a,8'h1a,8'h1a,8'h1a,8'h1a,8'h1a,8'h1a,8'h1a,8'h1a,8'h1a,8'h1a,8'h1a,8'h1a,8'h1a,8'h1a,8'h2b,8'h1a,8'h1a,8'h1a,8'h1a,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h1a,8'h1a,8'h1a,8'h1a,8'h1a,8'h1a,8'h1a,8'h1a,8'h1a,8'h21,8'h6,8'h6,8'h16,8'h3,8'h6,8'h2a,8'h1a,8'h1a,8'h1a,8'h2b,8'h1a,8'h1a,8'h9,8'h6,8'h9,8'h1a,8'h1a,8'h1a,8'h1a,8'h1a,8'h6,8'h6,8'h9,8'h2b,8'h2b,8'h1a,8'h1a,8'h1a,8'h22,8'h6,8'h9,8'h1a,8'h9,8'h6,8'h2a,8'h1a,8'h1a,8'h18,8'h22,8'h6,8'h21,8'h1a,8'h21,8'h6,8'h6,8'h1a,8'h1a,8'h1a,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h1a,8'h1a,8'h1a,8'h1a,8'h22,8'h6,8'h3,8'h2b,8'h1a,8'h2b,8'h1a,8'h3,8'h6,8'h9,8'h1a,8'h1a,8'h1a,8'h1a,8'h1a,8'h1a,8'h1a,8'h1a,8'h1a,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h1a,8'h1a,8'h1a,8'h1a,8'h1a,8'h2b,8'ha,8'h6,8'h22,8'h1a,8'h16,8'h6,8'h6,8'h2a,8'h1a,8'h1a,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h1a,8'h2b,8'h21,8'h6,8'h6,8'h1a,8'h1a,8'h1a,8'h1a,8'h1a,8'h1a,8'h1a,8'h1a,8'h16,8'h6,8'h6,8'h1b,8'h1a,8'h1a,8'h1a,8'h1a,8'h2b,8'h2b,8'h1a,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h1a,8'h1a,8'h1a,8'h16,8'h22,8'h1b,8'h1a,8'h1a,8'h1a,8'h6,8'h6,8'h9,8'h1a,8'h1a,8'h9,8'h6,8'h9,8'h16,8'h1a,8'h1a,8'h1a,8'h1a,8'h2,8'h6,8'h9,8'h1a,8'h1a,8'h1a,8'h1a,8'h1a,8'h22,8'h6,8'h21,8'h2b,8'h2b,8'h2b,8'h1a,8'h1a,8'h22,8'h6,8'h21,8'h2b,8'h16,8'h6,8'h6,8'h21,8'h1a,8'ha,8'h6,8'h6,8'h1a,8'h1a,8'h21,8'h6,8'h6,8'h1a,8'h1a,8'h1a,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h1a,8'h1a,8'h1a,8'h16,8'h21,8'h6,8'h6,8'h3,8'h2b,8'h2b,8'h9,8'h6,8'h6,8'h1b,8'h1a,8'h1a,8'h1a,8'h1a,8'h1a,8'h1a,8'h1a,8'h1a,8'h1a,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h1a,8'h1a,8'h1a,8'h2b,8'h3,8'h6,8'h9,8'h1a,8'h1a,8'h1b,8'h6,8'h6,8'h21,8'h1a,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h1a,8'h1a,8'h16,8'h6,8'h6,8'h1b,8'h1a,8'h1a,8'h21,8'h6,8'h2a,8'h1a,8'h1a,8'h16,8'h6,8'h6,8'h1b,8'h1a,8'h1a,8'h1a,8'h1a,8'h2b,8'h2b,8'h1a,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h1a,8'h1a,8'h1b,8'h6,8'h6,8'h6,8'h6,8'h6,8'h6,8'h21,8'h1a,8'h1a,8'h1a,8'h2b,8'h3,8'h6,8'h6,8'h6,8'h6,8'h6,8'h21,8'h9,8'h6,8'h9,8'h1a,8'h6,8'h6,8'h6,8'h6,8'h6,8'h9,8'h1a,8'h1b,8'h6,8'h6,8'h6,8'h6,8'h6,8'h9,8'h2b,8'h1a,8'h1a,8'h16,8'h6,8'h6,8'h6,8'h6,8'h22,8'h1a,8'h1a,8'h2b,8'h21,8'h6,8'h6,8'h1a,8'h2b,8'h1a,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h1a,8'h1a,8'h1a,8'h1a,8'h1a,8'h1a,8'h6,8'h6,8'h6,8'h6,8'h6,8'h9,8'h2b,8'h2b,8'h1a,8'h1a,8'h1a,8'h1a,8'h1a,8'h1a,8'h1a,8'h1a,8'h1a,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h1a,8'h2b,8'h1a,8'h1a,8'h2b,8'h1a,8'h3,8'h6,8'h22,8'h1a,8'h1a,8'h1a,8'h21,8'h6,8'h6,8'h21,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h1a,8'h1a,8'h16,8'h6,8'h6,8'h21,8'h1a,8'h1a,8'h9,8'h6,8'h6,8'h1a,8'h1a,8'h21,8'h6,8'h2a,8'h1a,8'h1a,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h1a,8'h2b,8'h1a,8'h2b,8'h1a,8'h1a,8'h1a,8'h1a,8'h1a,8'h2b,8'h1a,8'h1a,8'h2b,8'h2b,8'h2b,8'h1a,8'h1a,8'h2b,8'h2b,8'h2b,8'h1a,8'h1a,8'h1a,8'h1a,8'h1a,8'h1a,8'h2b,8'h1a,8'h1a,8'h2b,8'h2b,8'h1a,8'h2b,8'h1a,8'h2b,8'h1a,8'h1a,8'h2b,8'h2b,8'h1a,8'h1a,8'h1a,8'h1a,8'h1a,8'h1a,8'h1a,8'h2b,8'h1a,8'h1a,8'h1a,8'h1a,8'h1a,8'h1a,8'h1a,8'h1a,8'h1a,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h1a,8'h1a,8'h1a,8'h1a,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h1a,8'h1a,8'h1a,8'h2b,8'h1a,8'h1a,8'h1a,8'h1a,8'h1a,8'h1a,8'h1a,8'h1a,8'h1a,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h1a,8'h1a,8'h1a,8'h2b,8'h1a,8'h1a,8'h2b,8'h1a,8'h1a,8'h1a,8'h2b,8'h1a,8'h2b,8'h1a,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h1a,8'h1a,8'h18,8'h7,8'h6,8'h21,8'h1a,8'h16,8'h6,8'h6,8'h6,8'h1a,8'h1a,8'ha,8'h6,8'h2a,8'h1a,8'h2b,8'h1a,8'h1a,8'h2b,8'h1a,8'h1a,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h1a,8'h1a,8'h2b,8'h1a,8'h2b,8'h1a,8'h2b,8'h2b,8'h1a,8'h2b,8'h2b,8'h1a,8'h1a,8'h1a,8'h1a,8'h1a,8'h1a,8'h2b,8'h2b,8'h1a,8'h2b,8'h1a,8'h1a,8'h1a,8'h2b,8'h2b,8'h2b,8'h2b,8'h1a,8'h2b,8'h1a,8'h1a,8'h1a,8'h2b,8'h2b,8'h1a,8'h1a,8'h2b,8'h1a,8'h1a,8'h1a,8'h1a,8'h1a,8'h1a,8'h1a,8'h2b,8'h1a,8'h2b,8'h1a,8'h2b,8'h1a,8'h1a,8'h2b,8'h1a,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h1a,8'h1a,8'h1a,8'h1a,8'h2b,8'h1a,8'h2b,8'h1a,8'h1a,8'h1a,8'h1a,8'h1a,8'h2b,8'h1a,8'h1a,8'h1a,8'h1a,8'h1a,8'h1a,8'h1a,8'h1a,8'h1a,8'h1a,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h1a,8'h1a,8'h2b,8'h2b,8'h2b,8'h1a,8'h1a,8'h1a,8'h1a,8'h2b,8'h1a,8'h1a,8'h1a,8'h1a,8'h2b,8'h1a,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h1a,8'h18,8'h9,8'h6,8'h2a,8'h1a,8'h1b,8'h6,8'h6,8'h6,8'h2,8'h1a,8'h9,8'h6,8'h2a,8'h1a,8'h2b,8'h1a,8'h1a,8'h2b,8'h1a,8'h1a,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h1a,8'h2b,8'h1a,8'h1a,8'h2b,8'h1a,8'h2b,8'h1a,8'h1a,8'h2b,8'h1a,8'h1a,8'h1a,8'h1a,8'h1a,8'h1a,8'h1a,8'h2b,8'h2b,8'h1a,8'h1a,8'h2b,8'h1a,8'h2b,8'h2b,8'h1a,8'h1a,8'h2b,8'h1a,8'h2b,8'h1a,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h1a,8'h2b,8'h1a,8'h1a,8'h1a,8'h2b,8'h2b,8'h1a,8'h1a,8'h2b,8'h1a,8'h2b,8'h2b,8'h1a,8'h2b,8'h1a,8'h1a,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h1a,8'h1a,8'h1a,8'h1a,8'h2b,8'h2b,8'h1a,8'h1a,8'h2b,8'h2b,8'h1a,8'h1a,8'h2b,8'h1a,8'h1a,8'h1a,8'h1a,8'h1a,8'h1a,8'h1a,8'h1a,8'h1a,8'h1a,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h1a,8'h1a,8'h2b,8'h2b,8'h1a,8'h1a,8'h2b,8'h1a,8'h1a,8'h1a,8'h2b,8'h1a,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h1a,8'h1a,8'h1a,8'h4,8'h6,8'h2a,8'h1a,8'h3,8'h6,8'h6,8'h6,8'h2a,8'h1a,8'h22,8'h6,8'h21,8'h1a,8'h2b,8'h2b,8'h1a,8'h2b,8'h2b,8'h1a,8'h1a,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h1a,8'h2b,8'h1a,8'h2b,8'h1a,8'h2b,8'h2b,8'h1a,8'h2b,8'h2b,8'h1a,8'h1a,8'h1a,8'h1a,8'h1a,8'h1a,8'h1a,8'h1a,8'h1a,8'h2b,8'h2b,8'h1a,8'h2b,8'h1a,8'h1a,8'h2b,8'h2b,8'h2b,8'h1a,8'h2b,8'h2b,8'h2b,8'h1a,8'h1a,8'h2b,8'h2b,8'h1a,8'h2b,8'h1a,8'h2b,8'h2b,8'h1a,8'h1a,8'h1a,8'h2b,8'h2b,8'h1a,8'h2b,8'h2b,8'h1a,8'h2b,8'h1a,8'h2b,8'h2b,8'h1a,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h1a,8'h1a,8'h1a,8'h1a,8'h1a,8'h1a,8'h2b,8'h2b,8'h1a,8'h1a,8'h1a,8'h1a,8'h2b,8'h2b,8'h1a,8'h1a,8'h1a,8'h1a,8'h1a,8'h1a,8'h1a,8'h1a,8'h1a,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h1a,8'h2b,8'h2b,8'h2b,8'h2b,8'h1a,8'h2b,8'h2b,8'h1a,8'h2b,8'h1a,8'h2b,8'h1a,8'h2b,8'h1a,8'h1a,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h1a,8'h1a,8'h1a,8'h1b,8'h6,8'h6,8'h16,8'h22,8'h6,8'h6,8'h6,8'h6,8'h6,8'h6,8'h6,8'h1b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h1a,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h1a,8'h1a,8'h1a,8'h2b,8'h2b,8'h1a,8'h1a,8'h1a,8'h1a,8'h1a,8'h1a,8'h1a,8'h2b,8'h2b,8'h2b,8'h1a,8'h1a,8'h1a,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h1a,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h1a,8'h1a,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h1a,8'h1a,8'h1a,8'h1a,8'h2b,8'h1a,8'h1a,8'h2b,8'h1a,8'h1a,8'h1a,8'h1a,8'h1a,8'h2b,8'h1a,8'h1a,8'h1a,8'h1a,8'h1a,8'h1a,8'h1a,8'h1a,8'h1a,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h1a,8'h1a,8'h2b,8'h2b,8'h1a,8'h2b,8'h2b,8'h2b,8'h2b,8'h1a,8'h2b,8'h2b,8'h1a,8'h1a,8'h1a,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h1a,8'h1a,8'h1a,8'h1a,8'h6,8'h6,8'h6,8'h6,8'h22,8'h1a,8'h3,8'h6,8'h6,8'h6,8'h6,8'h1a,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h1a,8'h1a,8'h1a,8'h1a,8'h2b,8'h2b,8'h2b,8'h2b,8'h1a,8'h1a,8'h1a,8'h1a,8'h1a,8'h1a,8'h1a,8'h1a,8'h1a,8'h1a,8'h1a,8'h1a,8'h1a,8'h2b,8'h2b,8'h2b,8'h1a,8'h1a,8'h1a,8'h2b,8'h2b,8'h1a,8'h1a,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h1a,8'h1a,8'h2b,8'h2b,8'h2b,8'h1a,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h1a,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h1a,8'h1a,8'h1a,8'h1a,8'h2b,8'h2b,8'h2b,8'h1a,8'h1a,8'h2b,8'h1a,8'h1a,8'h1a,8'h1a,8'h1a,8'h1a,8'h1a,8'h1a,8'h1a,8'h1a,8'h1a,8'h1a,8'h1a,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h1a,8'h1a,8'h1a,8'h1a,8'h1a,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h1a,8'h1a,8'h1a,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h1a,8'h1a,8'h1a,8'h1a,8'h6,8'h6,8'h6,8'h6,8'h3,8'h2b,8'h21,8'h6,8'h6,8'h6,8'h22,8'h1a,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h1a,8'h1a,8'h2b,8'h1a,8'h2b,8'h2b,8'h2b,8'h1a,8'h1a,8'h2b,8'h1a,8'h1a,8'h1a,8'h1a,8'h2b,8'h2b,8'h2b,8'h1a,8'h1a,8'h2b,8'h2b,8'h2b,8'h2b,8'h1a,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h1a,8'h1a,8'h2b,8'h2b,8'h1a,8'h1a,8'h2b,8'h1a,8'h2b,8'h2b,8'h2b,8'h2b,8'h1a,8'h2b,8'h1a,8'h1a,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h1a,8'h1a,8'h1a,8'h1a,8'h1a,8'h1a,8'h1a,8'h1a,8'h1a,8'h2b,8'h1a,8'h1a,8'h2b,8'h1a,8'h1a,8'h1a,8'h1a,8'h1a,8'h1a,8'h1a,8'h1a,8'h1a,8'h1a,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h1a,8'h2b,8'h2b,8'h2b,8'h1a,8'h2b,8'h1a,8'h1a,8'h1a,8'h1a,8'h1a,8'h1a,8'h1a,8'h1a,8'h1a,8'h1a,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h1a,8'h1a,8'h1a,8'h2b,8'h3,8'h6,8'h6,8'h6,8'h1b,8'h1a,8'h16,8'h22,8'h6,8'h6,8'h21,8'h1a,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h1a,8'h1a,8'h1a,8'h1a,8'h1a,8'h1a,8'h1a,8'h1a,8'h1a,8'h1a,8'h1a,8'h2b,8'h2b,8'h1a,8'h1a,8'h1a,8'h2b,8'h1a,8'h1a,8'h1a,8'h2b,8'h2b,8'h1a,8'h1a,8'h2b,8'h2b,8'h1a,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h1a,8'h1a,8'h1a,8'h2b,8'h1a,8'h2b,8'h1a,8'h1a,8'h2b,8'h2b,8'h2b,8'h2b,8'h1a,8'h1a,8'h2b,8'h1a,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h1a,8'h1a,8'h1a,8'h1a,8'h1a,8'h2b,8'h2b,8'h2b,8'h2b,8'h1a,8'h1a,8'h1a,8'h2b,8'h2b,8'h1a,8'h1a,8'h1a,8'h1a,8'h1a,8'h1a,8'h1a,8'h1a,8'h1a,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h1a,8'h1a,8'h1a,8'h1a,8'h1a,8'h1a,8'h1a,8'h1a,8'h1a,8'h1a,8'h1a,8'h1a,8'h2b,8'h1a,8'h2b,8'h1a,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h1a,8'h1a,8'h1a,8'h2b,8'h16,8'h6,8'h6,8'h22,8'h1a,8'h1a,8'h16,8'h6,8'h6,8'h6,8'h21,8'h1a,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h1a,8'h1a,8'h1a,8'h3,8'h6,8'h6,8'h6,8'h6,8'h6,8'h21,8'h1a,8'h1a,8'h1a,8'h1a,8'h1a,8'h2b,8'h1a,8'h1a,8'h2b,8'h2b,8'h2b,8'h1a,8'h1a,8'h1a,8'h2b,8'h2b,8'h2b,8'h1a,8'h1a,8'h2b,8'h2b,8'h2b,8'h1a,8'h2b,8'h2b,8'h2b,8'h2b,8'h1a,8'h1a,8'h1a,8'h1a,8'h1a,8'h2b,8'h1a,8'h2b,8'h1a,8'h1a,8'h2b,8'h2b,8'h2b,8'h2b,8'h1a,8'h1a,8'h1a,8'h1a,8'h2b,8'h1a,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h1a,8'h1a,8'h1a,8'h1a,8'h2b,8'h21,8'h6,8'h6,8'h6,8'h6,8'h6,8'h6,8'h1b,8'h2b,8'h1a,8'h1a,8'h1a,8'h1a,8'h1a,8'h1a,8'h1a,8'h1a,8'h1a,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h1a,8'h1a,8'h2b,8'h2b,8'h1a,8'h21,8'h6,8'h6,8'h1a,8'h1a,8'h1a,8'h1a,8'h2b,8'h1a,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h1a,8'h1a,8'h1a,8'h1a,8'h1a,8'h1a,8'h1a,8'h2b,8'h1a,8'h1a,8'h1a,8'h1a,8'h1a,8'h1a,8'h1a,8'h1a,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h1a,8'h1a,8'h1a,8'h1a,8'h9,8'h6,8'h3,8'h1a,8'h1b,8'h6,8'h6,8'h3,8'h1a,8'h1a,8'h1a,8'h1a,8'h1a,8'h1a,8'h1a,8'h1a,8'h1a,8'h2b,8'h1a,8'h1a,8'h2b,8'h2b,8'h1a,8'h2b,8'h1a,8'h1a,8'h2b,8'h1a,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h1a,8'h1a,8'h1a,8'h1a,8'h1a,8'h2b,8'h1a,8'h1a,8'h1a,8'h1a,8'h2b,8'h2b,8'h2b,8'h2b,8'h1a,8'h1a,8'h1a,8'h1a,8'h2b,8'h1a,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h1a,8'h1a,8'h1a,8'h1a,8'h1a,8'h21,8'h6,8'h9,8'h1a,8'h2b,8'h21,8'h6,8'h6,8'h3,8'h1a,8'h1a,8'h1a,8'h1a,8'h1a,8'h1a,8'h1a,8'h1a,8'h1a,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h1a,8'h1a,8'h1a,8'h1a,8'h1a,8'h21,8'h6,8'h6,8'h1a,8'h1a,8'h1a,8'h1a,8'h2b,8'h1a,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h1a,8'h1a,8'h1a,8'h1a,8'h1a,8'h2b,8'h2b,8'h1a,8'h1a,8'h1a,8'h1a,8'h1a,8'h2b,8'h2b,8'h1a,8'h1a,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h1a,8'h1a,8'h1a,8'h1a,8'h9,8'h6,8'h9,8'h1a,8'h1a,8'h4,8'h6,8'h2a,8'h1a,8'h1a,8'h1a,8'h1a,8'h2b,8'h1a,8'h1a,8'h2b,8'h1a,8'h1a,8'h1a,8'h1a,8'h2b,8'h1a,8'h2b,8'h2b,8'h1a,8'h1a,8'h2b,8'h2b,8'h1a,8'h2b,8'h2b,8'h2b,8'h1a,8'h1a,8'h1a,8'h1a,8'h1a,8'h1a,8'h1a,8'h2b,8'h1a,8'h1a,8'h1a,8'h1a,8'h2b,8'h1a,8'h1a,8'h2b,8'h1a,8'h1a,8'h1a,8'h1a,8'h2b,8'h1a,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h1a,8'h1a,8'h1a,8'h1a,8'h2b,8'h21,8'h6,8'h9,8'h1a,8'h2b,8'h1a,8'h3,8'h6,8'h22,8'h1a,8'h1a,8'h1a,8'h1a,8'h1a,8'h1a,8'h1a,8'h1a,8'h1a,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h1a,8'h1a,8'h2b,8'h2b,8'h1a,8'h21,8'h6,8'h6,8'h1a,8'h1a,8'h1a,8'h1a,8'h1a,8'h1a,8'h2b,8'h1a,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h1a,8'h2b,8'h1a,8'h1a,8'h2b,8'h2b,8'h1a,8'h1a,8'h1a,8'h1a,8'h1a,8'h1a,8'h1a,8'h2b,8'h1a,8'h1a,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h1a,8'h1a,8'h1a,8'h1a,8'h9,8'h6,8'h9,8'h1a,8'h1a,8'h21,8'h6,8'h6,8'h1a,8'h21,8'h6,8'h2a,8'h1a,8'h1a,8'h16,8'h6,8'h6,8'h1b,8'h1a,8'h4,8'h6,8'h6,8'h6,8'h6,8'h6,8'h2,8'h1a,8'h2b,8'h1a,8'h2b,8'h2b,8'h2b,8'h1a,8'h1a,8'h1a,8'h1a,8'h1a,8'h1a,8'h1a,8'h2b,8'h1a,8'h1a,8'h1a,8'h1a,8'h2b,8'h1a,8'h1a,8'h2b,8'h1a,8'h1a,8'h1a,8'h1a,8'h2b,8'h1a,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h1a,8'h1a,8'h1a,8'h1a,8'h1a,8'h21,8'h6,8'h22,8'h1a,8'h1a,8'h1a,8'h21,8'h6,8'h6,8'h1a,8'h1a,8'h1a,8'h1a,8'h1a,8'h1a,8'h1a,8'h1a,8'h1a,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h1a,8'h1a,8'h2b,8'h1a,8'h1a,8'h21,8'h6,8'h6,8'h1a,8'h1a,8'h1a,8'h1a,8'h1a,8'h1a,8'h2b,8'h1a,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h1a,8'h1a,8'h1a,8'h1a,8'h1a,8'h2b,8'h2b,8'h1a,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h1a,8'h1a,8'h2b,8'h1a,8'h1a,8'h1a,8'h2b,8'h1a,8'h1a,8'h1a,8'h1a,8'h2b,8'h1a,8'h1a,8'h1a,8'h2b,8'h2b,8'h1a,8'h1a,8'h2b,8'h1a,8'h2b,8'h2b,8'h1a,8'h1a,8'h1a,8'h1a,8'h1a,8'h1a,8'h1a,8'h1a,8'h2b,8'h2b,8'h2b,8'h1a,8'h1a,8'h2b,8'h1a,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h1a,8'h1a,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h1a,8'h2b,8'h1a,8'h1a,8'h1a,8'h1a,8'h2b,8'h1a,8'h1a,8'h16,8'ha,8'h6,8'h9,8'h1a,8'h1a,8'ha,8'h6,8'h2a,8'h1a,8'h21,8'h6,8'h2a,8'h1a,8'h1a,8'h16,8'h6,8'h6,8'h1b,8'h1a,8'h21,8'h6,8'h2a,8'h1a,8'h1a,8'h9,8'h6,8'h2a,8'h1a,8'h2b,8'h1a,8'h1a,8'h2b,8'h1a,8'h1a,8'h1a,8'h1a,8'h2b,8'h1a,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h1a,8'h1a,8'h1a,8'h1a,8'h1a,8'h21,8'h6,8'h22,8'h1a,8'h1a,8'h1a,8'h3,8'h6,8'h6,8'h1a,8'h1a,8'h1a,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h1a,8'h1a,8'h1a,8'h1a,8'h1a,8'h21,8'h6,8'h6,8'h1a,8'h1a,8'h1a,8'h1a,8'h1a,8'h1a,8'h1a,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h1a,8'h1a,8'h1a,8'h1a,8'h1a,8'h1a,8'h1a,8'h1a,8'h1a,8'h1a,8'h1a,8'h1a,8'h1a,8'h1a,8'h1a,8'h1a,8'h2b,8'h2b,8'h1a,8'h2b,8'h1a,8'h1a,8'h1a,8'h2b,8'h2b,8'h1a,8'h1a,8'h1a,8'h2b,8'h2b,8'h1a,8'h1a,8'h1a,8'h1a,8'h2b,8'h1a,8'h1a,8'h2b,8'h1a,8'h1a,8'h1a,8'h1a,8'h1a,8'h1a,8'h1a,8'h2b,8'h1a,8'h1a,8'h1a,8'h2b,8'h1a,8'h1a,8'h1a,8'h1a,8'h1a,8'h2b,8'h1a,8'h1a,8'h2b,8'h1a,8'h1a,8'h1a,8'h1a,8'h1a,8'h1a,8'h2b,8'h1a,8'h2b,8'h1a,8'h1a,8'h1a,8'h1a,8'h1a,8'h1a,8'h1a,8'h1a,8'h1a,8'h2b,8'h1a,8'h1a,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h1a,8'h1a,8'h1a,8'h1a,8'h1a,8'h1a,8'h1a,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h1a,8'h2b,8'h1a,8'h1a,8'h1a,8'h1a,8'h1a,8'h2b,8'h1a,8'h1a,8'h1a,8'h1a,8'h2b,8'h1a,8'h1a,8'h1a,8'h2b,8'h2b,8'h1a,8'h1a,8'h2b,8'h1a,8'h2b,8'h1a,8'h1a,8'h1a,8'h1a,8'h1a,8'h1a,8'h1a,8'h1a,8'h1a,8'h2b,8'h1a,8'h2b,8'h2b,8'h2b,8'h2b,8'h1a,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h1a,8'h1a,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h1a,8'h2b,8'h1a,8'h1a,8'h1a,8'h1a,8'h2b,8'h1a,8'h1a,8'h1a,8'h9,8'h6,8'h9,8'h1a,8'h16,8'h6,8'h6,8'h3,8'h1a,8'h21,8'h6,8'h2a,8'h1a,8'h1a,8'h16,8'h6,8'h6,8'h1b,8'h1a,8'h21,8'h6,8'h2a,8'h1a,8'h1a,8'h21,8'h6,8'h6,8'h1a,8'h1a,8'h1a,8'h1a,8'h2b,8'h1a,8'h1a,8'h1a,8'h1a,8'h2b,8'h1a,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h1a,8'h1a,8'h1a,8'h1a,8'h1a,8'h21,8'h6,8'h22,8'h1a,8'h1a,8'h21,8'h6,8'h6,8'h3,8'h2b,8'h2b,8'h2b,8'h1a,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h1a,8'h1a,8'h1a,8'h1a,8'h1a,8'h21,8'h6,8'h6,8'h1a,8'h1a,8'h1a,8'h1a,8'h1a,8'h1a,8'h1a,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h1a,8'h1a,8'h3,8'h6,8'h6,8'h6,8'h6,8'h6,8'h1b,8'h1b,8'h1a,8'h1a,8'h2b,8'h1a,8'h1a,8'h1a,8'h2b,8'h2b,8'h2b,8'h2b,8'h1a,8'h1a,8'h1a,8'h1a,8'h1a,8'h2b,8'h1a,8'h1a,8'h1a,8'h2b,8'h1a,8'h1a,8'h1a,8'h2b,8'h1a,8'h1a,8'h2b,8'h1a,8'h1a,8'h1a,8'h2b,8'h2b,8'h1a,8'h1a,8'h1a,8'h2b,8'h1a,8'h1a,8'h2b,8'h1a,8'h1a,8'h1a,8'h21,8'h6,8'h6,8'h6,8'h6,8'h6,8'h6,8'h21,8'h1a,8'h1a,8'h1a,8'h1a,8'h1a,8'h2b,8'h1a,8'h2b,8'h1a,8'h2b,8'h1a,8'h1a,8'h2b,8'h1a,8'h1a,8'h1a,8'h1a,8'h1a,8'h1a,8'h1a,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h1a,8'h1a,8'h1a,8'h1a,8'h2b,8'h2b,8'h2b,8'h1a,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h1a,8'h2b,8'h2b,8'h2b,8'h1a,8'h1a,8'h1a,8'h1a,8'h1a,8'h1a,8'h1a,8'h1a,8'h1a,8'h1a,8'h1a,8'h1a,8'h2b,8'h2b,8'h1a,8'h1a,8'h2b,8'h1a,8'h2b,8'h1a,8'h1a,8'h2b,8'h1a,8'h1a,8'h1a,8'h1a,8'h1a,8'h1a,8'h2b,8'h1a,8'h1a,8'h1a,8'h1a,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h1a,8'h2b,8'h1a,8'h1a,8'h1a,8'h1a,8'h2b,8'h1a,8'h1a,8'h1a,8'h9,8'h6,8'h6,8'h6,8'h6,8'h6,8'h21,8'h1a,8'h1a,8'h21,8'h6,8'h2a,8'h1a,8'h1a,8'h16,8'h6,8'h6,8'h1b,8'h1a,8'h21,8'h6,8'h2a,8'h1a,8'h1a,8'h16,8'h6,8'h6,8'h1b,8'h1a,8'h1a,8'h1a,8'h2b,8'h1a,8'h1a,8'h1a,8'h1a,8'h2b,8'h1a,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h1a,8'h1a,8'h1a,8'h1a,8'h21,8'h6,8'h6,8'h6,8'h6,8'h6,8'h6,8'h21,8'h2b,8'h2b,8'h1a,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h1a,8'h1a,8'h1a,8'h1a,8'h1a,8'h21,8'h6,8'h6,8'h1a,8'h1a,8'h1a,8'h1a,8'h1a,8'h1a,8'h1a,8'h1a,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h1a,8'h9,8'h6,8'h22,8'h1a,8'h1a,8'h1a,8'h21,8'h1b,8'h1a,8'h1a,8'h1a,8'h1a,8'h1a,8'h1a,8'h1a,8'h1a,8'h1a,8'h1a,8'h1a,8'h1a,8'h1a,8'h1a,8'h2b,8'h2b,8'h1a,8'h2b,8'h2b,8'h1a,8'h1a,8'h1a,8'h1a,8'h1a,8'h2b,8'h1a,8'h2b,8'h2b,8'h2b,8'h1a,8'h1a,8'h1a,8'h2b,8'h1a,8'h1a,8'h1a,8'h2b,8'h1a,8'h1a,8'h2b,8'h1a,8'h1a,8'h1a,8'h21,8'h6,8'h6,8'h1a,8'h1a,8'h1a,8'h6,8'h6,8'h22,8'h1a,8'h1a,8'h1a,8'h2b,8'h2b,8'h1a,8'h1a,8'h2b,8'h2b,8'h1a,8'h2b,8'h1a,8'h1a,8'h2b,8'h1a,8'h1a,8'h1a,8'h1a,8'h1a,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h1a,8'h1a,8'h1a,8'h2b,8'h2b,8'h1a,8'h2b,8'h1a,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h1a,8'h2b,8'h1a,8'h1a,8'h1a,8'h2b,8'h2b,8'h1a,8'h1a,8'h1a,8'h1a,8'h2b,8'h1a,8'h1a,8'h1a,8'h2b,8'h2b,8'h1a,8'h1a,8'h2b,8'h1a,8'h2b,8'h1a,8'h1a,8'h1a,8'h1a,8'h1a,8'h1a,8'h1a,8'h1a,8'h1a,8'h2b,8'h2b,8'h2b,8'h2b,8'h1a,8'h2b,8'h2b,8'h1a,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h1a,8'h2b,8'h1a,8'h1a,8'h1a,8'h1a,8'h2b,8'h1a,8'h1a,8'h1a,8'h9,8'h6,8'h2,8'h21,8'h6,8'h6,8'h21,8'h1a,8'h1a,8'h21,8'h6,8'h22,8'h1a,8'h1a,8'h16,8'h6,8'h6,8'h1b,8'h1a,8'h21,8'h6,8'h2a,8'h1a,8'h1a,8'h16,8'h6,8'h6,8'h1b,8'h2b,8'h1a,8'h1a,8'h2b,8'h1a,8'h1a,8'h1a,8'h1a,8'h2b,8'h1a,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h1a,8'h1a,8'h1a,8'h1a,8'h21,8'h6,8'h9,8'h1a,8'h1a,8'h2b,8'h2b,8'h2b,8'h1a,8'h1a,8'h2b,8'h2b,8'h1a,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h1a,8'h1a,8'h1a,8'h1a,8'h1a,8'h21,8'h6,8'h6,8'h1a,8'h1a,8'h1a,8'h1a,8'h1a,8'h2b,8'h2b,8'h1a,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h16,8'h6,8'h6,8'h1b,8'h2b,8'h1a,8'h1a,8'h1a,8'h1a,8'h1a,8'h1a,8'h1a,8'h1a,8'h1a,8'h1a,8'h1a,8'h2b,8'h1a,8'h2b,8'h1a,8'h1a,8'h1a,8'h1a,8'h1a,8'h1a,8'h2b,8'h1a,8'h1a,8'h1a,8'h1a,8'h1a,8'h1a,8'h1a,8'h2b,8'h1a,8'h1a,8'h1a,8'h2b,8'h1a,8'h1a,8'h2b,8'h2b,8'h1a,8'h1a,8'h2b,8'h1a,8'h1a,8'h1a,8'h2b,8'h1a,8'h1a,8'h1a,8'h21,8'h6,8'h22,8'h1a,8'h2b,8'h1a,8'h1b,8'h6,8'h6,8'h1b,8'h1a,8'h16,8'h1a,8'h1a,8'h1a,8'h1a,8'h1a,8'h1a,8'h1a,8'h1a,8'h1a,8'h1a,8'h1a,8'h1a,8'h1a,8'h1a,8'h2b,8'h1a,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h1a,8'h1a,8'h1a,8'h1a,8'h1a,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h1a,8'h1a,8'h1a,8'h1a,8'h1a,8'h1a,8'h1a,8'h1a,8'h1a,8'h2b,8'h1a,8'h2b,8'h2b,8'h2b,8'h2b,8'h1a,8'h1a,8'h2b,8'h1a,8'h2b,8'h1a,8'h1a,8'h1a,8'h1a,8'h1a,8'h1a,8'h1a,8'h1a,8'h1a,8'h1a,8'h1a,8'h2b,8'h2b,8'h2b,8'h1a,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h1a,8'h2b,8'h1a,8'h1a,8'h1a,8'h1a,8'h2b,8'h1a,8'h1a,8'h1a,8'ha,8'h6,8'h9,8'h1a,8'h21,8'h6,8'h6,8'h1b,8'h1a,8'h1b,8'h6,8'h6,8'h1a,8'h1a,8'h16,8'h6,8'h6,8'h1b,8'h1a,8'h21,8'h6,8'h2a,8'h1a,8'h1a,8'h16,8'h6,8'h6,8'h1b,8'h2b,8'h1a,8'h1a,8'h2b,8'h1a,8'h1a,8'h1a,8'h1a,8'h2b,8'h1a,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h1a,8'h1a,8'h1a,8'h1a,8'h21,8'h6,8'h9,8'h1a,8'h1a,8'h1a,8'h2b,8'h2b,8'h1a,8'h2b,8'h2b,8'h1a,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h1a,8'h1a,8'h1a,8'h1a,8'h1a,8'h21,8'h6,8'h6,8'h1a,8'h1a,8'h1a,8'h1a,8'h1a,8'h1a,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h1a,8'h22,8'h6,8'h22,8'h1a,8'h1a,8'h1a,8'h2b,8'h1a,8'h1a,8'h21,8'h6,8'h6,8'h6,8'h6,8'h6,8'h6,8'h1a,8'h1a,8'h1a,8'h16,8'h6,8'h6,8'h6,8'h6,8'h6,8'h1b,8'h1a,8'h1a,8'h1a,8'h1a,8'h3,8'h6,8'h6,8'h6,8'h6,8'h6,8'h1b,8'h1a,8'h1a,8'h6,8'h6,8'h6,8'h6,8'h6,8'h1b,8'h1a,8'h1a,8'h1a,8'h1a,8'h1a,8'h1a,8'h21,8'h6,8'h6,8'h1a,8'h2b,8'h1a,8'h1b,8'h6,8'h6,8'h1b,8'h1a,8'h16,8'h6,8'h6,8'h6,8'h6,8'h6,8'h1b,8'h1a,8'h1a,8'h21,8'h6,8'h6,8'h6,8'h6,8'h6,8'h3,8'h1a,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h1a,8'h1a,8'h1a,8'h1a,8'h1a,8'h2b,8'h2b,8'h2b,8'h2b,8'h1a,8'h1a,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h1a,8'h2b,8'h1a,8'h4,8'h6,8'h6,8'h6,8'h6,8'h22,8'h21,8'h2b,8'h1a,8'h2b,8'h1a,8'h2b,8'h2b,8'h1a,8'h1a,8'h2b,8'h1a,8'h2b,8'h1a,8'h1a,8'h1a,8'h1a,8'h1a,8'h1a,8'h1a,8'h1a,8'h1a,8'h2b,8'h2b,8'h1a,8'h1a,8'h2b,8'h1a,8'h1a,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h1a,8'h1a,8'h1a,8'h1a,8'h2b,8'h1a,8'h1a,8'h1a,8'h9,8'h6,8'h9,8'h1a,8'h1a,8'h9,8'h6,8'h22,8'h1a,8'h1a,8'h6,8'h6,8'h22,8'h1a,8'h16,8'h6,8'h6,8'h1b,8'h1a,8'h21,8'h6,8'h22,8'h1a,8'h1a,8'h16,8'h6,8'h6,8'h1b,8'h1a,8'h1a,8'h1a,8'h2b,8'h1a,8'h1a,8'h1a,8'h1a,8'h2b,8'h1a,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h1a,8'h1a,8'h1a,8'h1a,8'h21,8'h6,8'h22,8'h1a,8'h1a,8'h2b,8'h1a,8'h1a,8'h2b,8'h2b,8'h2b,8'h1a,8'h1a,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h1a,8'h1a,8'h1a,8'h1a,8'h1a,8'h21,8'h6,8'h6,8'h1a,8'h1a,8'h1a,8'h1a,8'h1a,8'h2b,8'h2b,8'h1a,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h1a,8'h21,8'h6,8'h6,8'h6,8'h6,8'h6,8'h1b,8'h1a,8'h1a,8'h21,8'h6,8'h2a,8'h1a,8'h1a,8'h9,8'h6,8'h6,8'h1a,8'h1a,8'h18,8'h1a,8'h2b,8'h1a,8'h3,8'h6,8'h6,8'h1a,8'h1a,8'h1a,8'h6,8'h6,8'h2,8'h1a,8'h16,8'h1a,8'h1a,8'h2b,8'h1a,8'h6,8'h6,8'h21,8'h2b,8'h21,8'h6,8'h6,8'h1b,8'h1a,8'h1a,8'h1a,8'h1a,8'h1a,8'h21,8'h6,8'h6,8'h1a,8'h1a,8'h1a,8'h22,8'h6,8'h2a,8'h1a,8'h1a,8'h1a,8'h1a,8'h1a,8'h1a,8'h3,8'h6,8'h6,8'h1a,8'h1a,8'h21,8'h6,8'h6,8'h1b,8'h2b,8'h1a,8'h1a,8'h1a,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h1a,8'h1a,8'h1a,8'h1a,8'h2b,8'h1a,8'h2b,8'h1a,8'h2b,8'h2b,8'h1a,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h1a,8'h1a,8'h2b,8'h2b,8'h1a,8'h9,8'h6,8'h9,8'h1a,8'h1a,8'h1b,8'h21,8'h1b,8'h1a,8'h1a,8'h2b,8'h2b,8'h2b,8'h2b,8'h1a,8'h1a,8'h2b,8'h2b,8'h2b,8'h1a,8'h21,8'h6,8'h6,8'h6,8'h6,8'h6,8'h6,8'h21,8'h1a,8'h2b,8'h2b,8'h1a,8'h2b,8'h2b,8'h1a,8'h1a,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h1a,8'h1a,8'h1a,8'h1a,8'h2b,8'h1a,8'h1a,8'h1a,8'h9,8'h6,8'h9,8'h1a,8'h1a,8'h1b,8'h6,8'h6,8'h21,8'h2b,8'h1a,8'h3,8'h6,8'h6,8'h6,8'h6,8'h3,8'h1a,8'h1a,8'h21,8'h6,8'h22,8'h1a,8'h1a,8'h1a,8'h6,8'h6,8'h1b,8'h2b,8'h1a,8'h1a,8'h2b,8'h1a,8'h1a,8'h1a,8'h1a,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h1a,8'h1a,8'h1a,8'h1a,8'h21,8'h6,8'h9,8'h1a,8'h1a,8'h2b,8'h1a,8'h2b,8'h2b,8'h1a,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h1a,8'h1a,8'h1a,8'h1a,8'h1a,8'h21,8'h6,8'h6,8'h6,8'h6,8'h6,8'h6,8'h6,8'h3,8'h1a,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h1a,8'h1a,8'h16,8'h6,8'h6,8'h6,8'h6,8'h6,8'h3,8'h1a,8'h21,8'h6,8'h2a,8'h1a,8'h1a,8'h1a,8'h22,8'h6,8'h21,8'h1a,8'h1a,8'h1a,8'h1a,8'h1a,8'h16,8'h6,8'h6,8'h1a,8'h1a,8'h21,8'h6,8'h22,8'h1a,8'h1a,8'h1a,8'h1a,8'h1a,8'h1a,8'h4,8'h6,8'h9,8'h2b,8'h1a,8'h1a,8'h9,8'h6,8'h21,8'h1a,8'h1a,8'h1a,8'h2b,8'h1a,8'h1,8'h6,8'h6,8'h6,8'h6,8'h6,8'h6,8'h22,8'h1a,8'h1a,8'h1a,8'h1a,8'h1a,8'h2b,8'h1a,8'h16,8'h6,8'h6,8'h1b,8'h1a,8'h21,8'h6,8'h6,8'h1a,8'h1a,8'h1a,8'h1a,8'h1a,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h1a,8'h1a,8'h1a,8'h1a,8'h1a,8'h1b,8'h6,8'h6,8'h6,8'h1b,8'h1a,8'h2b,8'h1a,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h1a,8'h1a,8'h2b,8'h1a,8'h2b,8'h16,8'h6,8'h6,8'h21,8'h2b,8'h1a,8'h1a,8'h1a,8'h1a,8'h1a,8'h1a,8'h2b,8'h2b,8'h2b,8'h2b,8'h1a,8'h1a,8'h2b,8'h2b,8'h1a,8'h1a,8'h21,8'h6,8'h6,8'h1a,8'h1a,8'h1a,8'h6,8'h6,8'h6,8'h1b,8'h2b,8'h1a,8'h1a,8'h2b,8'h2b,8'h1a,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h1a,8'h1a,8'h2b,8'h1a,8'h2b,8'h1a,8'h1a,8'h2b,8'h1a,8'h1a,8'h1a,8'h1a,8'h1a,8'h1a,8'h1a,8'h1a,8'h1a,8'h2b,8'h1a,8'h1a,8'h1a,8'h1a,8'h1a,8'h1a,8'h1a,8'h1a,8'h1a,8'h1a,8'h1a,8'h1a,8'h1a,8'h1a,8'h1a,8'h1a,8'h1a,8'h1a,8'h1a,8'h1a,8'h1a,8'h1a,8'h1a,8'h1a,8'h1a,8'h1a,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h1a,8'h1a,8'h1a,8'h1a,8'h1a,8'h2b,8'h1a,8'h1a,8'h1a,8'h1a,8'h2b,8'h1a,8'h2b,8'h2b,8'h1a,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h1a,8'h1a,8'h1a,8'h1a,8'h1a,8'h2b,8'h1a,8'h2b,8'h1a,8'h1a,8'h1a,8'h1a,8'h1a,8'h2b,8'h2b,8'h1a,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h1a,8'h1a,8'h1a,8'h2b,8'h1a,8'h1a,8'h22,8'h6,8'h6,8'h1a,8'h0,8'h6,8'h2a,8'h1a,8'h1a,8'h1a,8'h9,8'h6,8'h2a,8'h1a,8'h1a,8'h22,8'h6,8'h6,8'h6,8'h6,8'h6,8'h1b,8'h1a,8'h9,8'h6,8'h2a,8'h1a,8'h1a,8'h1a,8'h1a,8'h2b,8'h1a,8'h22,8'h6,8'h6,8'h6,8'h6,8'h6,8'h6,8'h6,8'h9,8'h1a,8'h1a,8'h1a,8'h1a,8'h1a,8'h21,8'h6,8'h6,8'h1a,8'h2b,8'h1a,8'h21,8'h6,8'h6,8'h21,8'h1a,8'h18,8'h6,8'h6,8'h6,8'h6,8'h6,8'h6,8'h1a,8'h1a,8'h21,8'h6,8'h6,8'h1a,8'h1a,8'h1a,8'h1a,8'h1a,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h1a,8'h2b,8'h2b,8'h1a,8'h1a,8'h1a,8'h1a,8'h1a,8'h3,8'h6,8'h6,8'h6,8'h21,8'h2b,8'h2b,8'h1a,8'h1a,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h1a,8'h1a,8'h1a,8'h2b,8'h2b,8'h1a,8'h22,8'h6,8'h22,8'h2b,8'h1a,8'h1a,8'h1a,8'h1a,8'h1a,8'h1a,8'h2b,8'h1a,8'h1a,8'h2b,8'h1a,8'h1a,8'h2b,8'h2b,8'h1a,8'h1a,8'h21,8'h6,8'h6,8'h1a,8'h1a,8'h1a,8'h1a,8'h9,8'h6,8'h9,8'h1a,8'h1a,8'h1a,8'h2b,8'h1a,8'h1a,8'h1a,8'h1a,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h1a,8'h1a,8'h2b,8'h2b,8'h2b,8'h1a,8'h1a,8'h2b,8'h1a,8'h1a,8'h1a,8'h1a,8'h1a,8'h1a,8'h1a,8'h2b,8'h2b,8'h2b,8'h1a,8'h1a,8'h1a,8'h2b,8'h1a,8'h1a,8'h1a,8'h1a,8'h2b,8'h1a,8'h1a,8'h1a,8'h1a,8'h1a,8'h1a,8'h1a,8'h1a,8'h1a,8'h2b,8'h2b,8'h1a,8'h1a,8'h1a,8'h1a,8'h1a,8'h1a,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h1a,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h1a,8'h1a,8'h1a,8'h1a,8'h2b,8'h2b,8'h1a,8'h1a,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h1a,8'h1a,8'h1a,8'h1a,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h1a,8'h1a,8'h1a,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h1a,8'h1a,8'h1a,8'h1a,8'h1a,8'h1a,8'h21,8'h6,8'h6,8'h1b,8'h21,8'h6,8'h22,8'h1a,8'h1a,8'h1a,8'h9,8'h6,8'h3,8'h1a,8'h6,8'h6,8'h2a,8'h1a,8'h16,8'h6,8'h6,8'h1b,8'h1a,8'h9,8'h6,8'h2a,8'h1a,8'h1a,8'h1a,8'h1a,8'h2b,8'h1a,8'h22,8'h6,8'h21,8'h2b,8'h1a,8'h2b,8'h2b,8'h1a,8'h1a,8'h1a,8'h1a,8'h1a,8'h1a,8'h1a,8'h21,8'h6,8'h6,8'h1a,8'h1a,8'h1a,8'h1a,8'h9,8'h6,8'h2,8'h16,8'h22,8'h6,8'h3,8'h1a,8'h16,8'h6,8'h6,8'h1b,8'h1a,8'h0,8'h6,8'h6,8'h1a,8'h2b,8'h1a,8'h1a,8'h1a,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h1a,8'h1a,8'h1a,8'h1a,8'h1a,8'h22,8'h6,8'h6,8'h6,8'h22,8'h1a,8'h1a,8'h1a,8'h1a,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h1a,8'h1a,8'h1a,8'h1a,8'h2b,8'h1a,8'h21,8'h6,8'h6,8'h6,8'h6,8'h6,8'h1b,8'h1a,8'h1a,8'h1a,8'h2b,8'h2b,8'h1a,8'h2b,8'h1a,8'h1a,8'h2b,8'h1a,8'h1a,8'h1a,8'h1,8'h6,8'h6,8'h1a,8'h1a,8'h1a,8'h1a,8'h16,8'h6,8'h6,8'h21,8'h1a,8'h1a,8'h2b,8'h1a,8'h1a,8'h1a,8'h1a,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h1a,8'h2b,8'h2b,8'h2b,8'h2b,8'h1a,8'h1a,8'h2b,8'h2b,8'h2b,8'h1a,8'h1a,8'h1a,8'h2b,8'h1a,8'h2b,8'h2b,8'h2b,8'h1a,8'h1a,8'h2b,8'h2b,8'h1a,8'h1a,8'h1a,8'h1a,8'h2b,8'h2b,8'h2b,8'h1a,8'h1a,8'h1a,8'h1a,8'h2b,8'h2b,8'h1a,8'h2b,8'h2b,8'h2b,8'h1a,8'h1a,8'h1a,8'h1a,8'h1a,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h1a,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h1a,8'h1a,8'h1a,8'h1a,8'h2b,8'h2b,8'h1a,8'h1a,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h1a,8'h1a,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h1a,8'h1a,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h1a,8'h1a,8'h1a,8'h2b,8'h1a,8'h1a,8'h21,8'h6,8'h6,8'h1a,8'h21,8'h6,8'h22,8'h1a,8'h2b,8'h1a,8'h22,8'h6,8'h3,8'h1a,8'h6,8'h6,8'h1b,8'h1a,8'h16,8'h6,8'h6,8'h1b,8'h1a,8'h3,8'h6,8'h22,8'h1a,8'h1a,8'h1a,8'h1a,8'h2b,8'h1a,8'h3,8'h6,8'h22,8'h1a,8'h2b,8'h1a,8'h2b,8'h1a,8'h1a,8'h1a,8'h1a,8'h1a,8'h1a,8'h1a,8'h21,8'h6,8'h6,8'h1a,8'h2b,8'h1a,8'h1a,8'hb,8'h6,8'h2a,8'h16,8'h7,8'h6,8'h21,8'h1a,8'h16,8'h6,8'h6,8'h1a,8'h1a,8'h21,8'h6,8'h6,8'h1a,8'h2b,8'h1a,8'h1a,8'h1a,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h1a,8'h2b,8'h1a,8'h1a,8'h1a,8'h1a,8'h21,8'h6,8'h6,8'h21,8'h6,8'h6,8'h1b,8'h1a,8'h1a,8'h1a,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h1a,8'h1a,8'h1a,8'h2b,8'h2b,8'h1a,8'h1a,8'h16,8'h6,8'h6,8'h6,8'h6,8'h6,8'h21,8'h1a,8'h1a,8'h2b,8'h2b,8'h1a,8'h2b,8'h1a,8'h1a,8'h2b,8'h1a,8'h1a,8'h1a,8'h21,8'h6,8'h6,8'h1a,8'h1a,8'h1a,8'h1a,8'h1a,8'h6,8'h6,8'h3,8'h1a,8'h1a,8'h1a,8'h1a,8'h1a,8'h1a,8'h1a,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h1a,8'h2b,8'h2b,8'h2b,8'h1a,8'h1a,8'h2b,8'h2b,8'h1a,8'h1a,8'h2b,8'h1a,8'h2b,8'h2b,8'h2b,8'h2b,8'h1a,8'h1a,8'h1a,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h1a,8'h1a,8'h1a,8'h1a,8'h1a,8'h1a,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h1a,8'h1a,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h1a,8'h1a,8'h1a,8'h1a,8'h2b,8'h2b,8'h1a,8'h1a,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h1a,8'h1a,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h1a,8'h1a,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h16,8'h22,8'h16,8'h2b,8'h1a,8'h1a,8'h6,8'h6,8'h2a,8'h1a,8'h21,8'h6,8'h6,8'h1a,8'h1a,8'h4,8'h6,8'h6,8'h1a,8'h1a,8'h7,8'h6,8'h21,8'h1a,8'h16,8'h6,8'h6,8'h1b,8'h2b,8'h1a,8'h22,8'h6,8'h9,8'h1a,8'h1a,8'h1a,8'h1a,8'h2b,8'h16,8'h6,8'h6,8'h2,8'h1a,8'h2b,8'h1a,8'h1a,8'h1a,8'h1a,8'h1a,8'h1a,8'h1a,8'h1a,8'h21,8'h6,8'h22,8'h1a,8'h2b,8'h16,8'h21,8'h6,8'h6,8'h1b,8'h1a,8'h6,8'h6,8'h21,8'h16,8'h16,8'h22,8'h6,8'h1b,8'h1a,8'h21,8'h6,8'h6,8'h1a,8'h1a,8'h1a,8'h2b,8'h1a,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h1a,8'h2b,8'h1a,8'h1a,8'h1a,8'h1a,8'h9,8'h6,8'h9,8'h2b,8'h6,8'h6,8'h21,8'h1a,8'h1a,8'h1a,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h1a,8'h1a,8'h1a,8'h1a,8'h2b,8'h1a,8'h1a,8'h1a,8'h1a,8'h1a,8'h1a,8'h6,8'h6,8'h6,8'h1a,8'h1a,8'h1a,8'h1a,8'h1a,8'h2b,8'h1a,8'h1a,8'h2b,8'h1a,8'h1a,8'h1a,8'h21,8'h6,8'h6,8'h1a,8'h1a,8'h1a,8'h1a,8'h18,8'h22,8'h6,8'h3,8'h1a,8'h1a,8'h1a,8'h1a,8'h1a,8'h1a,8'h1a,8'h1a,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h1a,8'h2b,8'h2b,8'h2b,8'h1a,8'h1a,8'h2b,8'h2b,8'h1a,8'h1a,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h1a,8'h1a,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h1a,8'h1a,8'h1a,8'h1a,8'h1a,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h1a,8'h1a,8'h2b,8'h2b,8'h2b,8'h1a,8'h2b,8'h2b,8'h2b,8'h1a,8'h1a,8'h1a,8'h2b,8'h2b,8'h1a,8'h1a,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h1a,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h1a,8'h1a,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h16,8'h6,8'h6,8'h6,8'h6,8'h6,8'h6,8'h3,8'h1a,8'h1a,8'h4,8'h6,8'h6,8'h6,8'h6,8'h6,8'h22,8'h1a,8'h1a,8'h1a,8'h16,8'h6,8'h6,8'h6,8'h6,8'h6,8'h6,8'h1a,8'h1a,8'h1a,8'h16,8'ha,8'h6,8'h6,8'h6,8'h6,8'h6,8'h21,8'h1a,8'h1a,8'h22,8'h6,8'h6,8'h6,8'h6,8'h6,8'h1a,8'h1a,8'h1a,8'h2b,8'h2b,8'h1a,8'h21,8'h6,8'h6,8'h6,8'h6,8'h6,8'h6,8'h6,8'h1a,8'h1a,8'h1a,8'h18,8'h6,8'h6,8'h6,8'h22,8'h6,8'h6,8'h1b,8'h1a,8'h21,8'h6,8'h6,8'h1a,8'h2b,8'h1a,8'h1a,8'h1a,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h1a,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h1a,8'h1a,8'h1a,8'h1a,8'h1a,8'h1a,8'h16,8'h6,8'h6,8'h21,8'h1a,8'h3,8'h6,8'h22,8'h1a,8'h1a,8'h1a,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h1a,8'h1a,8'h1a,8'h1a,8'h1a,8'h1a,8'h1a,8'h1a,8'h1a,8'h1a,8'h1a,8'h21,8'h6,8'h22,8'h1b,8'h1a,8'h1a,8'h1a,8'h1a,8'h2b,8'h1a,8'h1a,8'h2b,8'h1a,8'h1a,8'h1a,8'h0,8'h6,8'h6,8'h1a,8'h2b,8'h1a,8'h1a,8'h1a,8'h22,8'h6,8'h21,8'h1a,8'h1a,8'h1a,8'h1a,8'h1a,8'h1a,8'h1a,8'h1a,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h1a,8'h2b,8'h2b,8'h2b,8'h1a,8'h1a,8'h2b,8'h2b,8'h1a,8'h1a,8'h2b,8'h2b,8'h1a,8'h1a,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h1a,8'h1a,8'h1a,8'h1a,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h1a,8'h1a,8'h2b,8'h2b,8'h2b,8'h1a,8'h2b,8'h2b,8'h2b,8'h1a,8'h1a,8'h1a,8'h2b,8'h2b,8'h1a,8'h1a,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h1a,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h1a,8'h1a,8'h1a,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h1a,8'h1a,8'h1a,8'h1a,8'h1a,8'h1a,8'h2b,8'h2b,8'h1a,8'h1a,8'h21,8'h6,8'h22,8'h1a,8'h1a,8'h1a,8'h2b,8'h1a,8'h1a,8'h2b,8'h1a,8'h1a,8'h2b,8'h1a,8'h1a,8'h2b,8'h1a,8'h1a,8'h1a,8'h1a,8'h1a,8'h1a,8'h1a,8'h1a,8'h1a,8'h1a,8'h1a,8'h2b,8'h1a,8'h1a,8'h2b,8'h1a,8'h1a,8'h1a,8'h1a,8'h2b,8'h1a,8'h1a,8'h2b,8'h1a,8'h1a,8'h1a,8'h1a,8'h1a,8'h1a,8'h1a,8'h1a,8'h1a,8'h1a,8'h2b,8'h1a,8'h1a,8'h1a,8'h1a,8'h2b,8'h1a,8'h1a,8'h1a,8'h1a,8'h2b,8'h1a,8'h1a,8'h1a,8'h1a,8'h1a,8'h1a,8'h1a,8'h2b,8'h2b,8'h1a,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h1a,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h1a,8'h2b,8'h1a,8'h1a,8'h1a,8'h1a,8'h21,8'h6,8'h6,8'h1a,8'h1a,8'h1b,8'h6,8'h6,8'h1b,8'h1a,8'h1a,8'h1a,8'h2b,8'h2b,8'h2b,8'h2b,8'h1a,8'h1a,8'h1a,8'h1a,8'h1a,8'h1a,8'h1a,8'h1a,8'h1a,8'h1a,8'h1a,8'h21,8'h6,8'h6,8'h1a,8'h1a,8'h1a,8'h1a,8'h1a,8'h2b,8'h1a,8'h1a,8'h2b,8'h1a,8'h1a,8'h1a,8'h21,8'h6,8'h6,8'h1a,8'h2b,8'h1a,8'h1a,8'h21,8'h6,8'h6,8'h21,8'h1a,8'h1a,8'h1a,8'h1a,8'h1a,8'h1a,8'h1a,8'h1a,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h1a,8'h2b,8'h2b,8'h2b,8'h1a,8'h1a,8'h2b,8'h2b,8'h1a,8'h1a,8'h2b,8'h2b,8'h1a,8'h1a,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h1a,8'h1a,8'h1a,8'h1a,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h1a,8'h1a,8'h2b,8'h2b,8'h2b,8'h1a,8'h2b,8'h2b,8'h2b,8'h1a,8'h1a,8'h1a,8'h2b,8'h2b,8'h1a,8'h1a,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h1a,8'h1a,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h1a,8'h1a,8'h1a,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h1a,8'h1a,8'h1a,8'h1a,8'h1a,8'h2b,8'h2b,8'h2b,8'h1a,8'h1a,8'h21,8'h6,8'h9,8'h1a,8'h2b,8'h1a,8'h1a,8'h2b,8'h2b,8'h2b,8'h1a,8'h1a,8'h1a,8'h2b,8'h2b,8'h1a,8'h1a,8'h2b,8'h1a,8'h1a,8'h1a,8'h1a,8'h1a,8'h2b,8'h1a,8'h2b,8'h2b,8'h2b,8'h1a,8'h1a,8'h1a,8'h2b,8'h1a,8'h1a,8'h2b,8'h1a,8'h1a,8'h1a,8'h1a,8'h1a,8'h1a,8'h1a,8'h1a,8'h2b,8'h1a,8'h1a,8'h2b,8'h1a,8'h2b,8'h1a,8'h1a,8'h1a,8'h1a,8'h1a,8'h1a,8'h2b,8'h1a,8'h1a,8'h1a,8'h2b,8'h1a,8'h2b,8'h1a,8'h1a,8'h2b,8'h1a,8'h2b,8'h1a,8'h1a,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h1a,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h1a,8'h2b,8'h1a,8'h1a,8'h1a,8'h1a,8'h9,8'h6,8'h6,8'h6,8'h6,8'h6,8'h6,8'h6,8'h3,8'h1a,8'h1a,8'h1a,8'h2b,8'h2b,8'h2b,8'h2b,8'h1a,8'h1a,8'h1a,8'h1a,8'h1a,8'h1a,8'h6,8'h16,8'h1a,8'h1a,8'h1a,8'h6,8'h6,8'h2a,8'h1a,8'h1a,8'h1a,8'h1a,8'h1a,8'h2b,8'h1a,8'h1a,8'h2b,8'h1a,8'h1a,8'h1a,8'h0,8'h6,8'h2a,8'h1a,8'h1a,8'h1a,8'h16,8'h23,8'h6,8'h2a,8'h1a,8'h1a,8'h1a,8'h1a,8'h1a,8'h1a,8'h1a,8'h1a,8'h1a,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h1a,8'h1a,8'h1a,8'h1a,8'h1a,8'h1a,8'h2b,8'h2b,8'h1a,8'h1a,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h1a,8'h1a,8'h1a,8'h1a,8'h1a,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h1a,8'h1a,8'h2b,8'h2b,8'h2b,8'h1a,8'h2b,8'h2b,8'h2b,8'h1a,8'h1a,8'h1a,8'h2b,8'h2b,8'h1a,8'h1a,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h1a,8'h1a,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h1a,8'h1a,8'h1a,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h1a,8'h1a,8'h1a,8'h1a,8'h1a,8'h1a,8'h1a,8'h1a,8'h2b,8'h1a,8'h1a,8'h1a,8'h1a,8'h1a,8'h1a,8'h2b,8'h2b,8'h2b,8'h1a,8'h1a,8'h1a,8'h1a,8'h1a,8'h2b,8'h2b,8'h1a,8'h2b,8'h2b,8'h1a,8'h2b,8'h1a,8'h1a,8'h1a,8'h1a,8'h1a,8'h2b,8'h2b,8'h1a,8'h1a,8'h1a,8'h2b,8'h1a,8'h1a,8'h1a,8'h1a,8'h2b,8'h1a,8'h1a,8'h1a,8'h1a,8'h1a,8'h1a,8'h1a,8'h1a,8'h1a,8'h1a,8'h2b,8'h1a,8'h1a,8'h2b,8'h1a,8'h1a,8'h1a,8'h1a,8'h2b,8'h1a,8'h1a,8'h1a,8'h1a,8'h1a,8'h1a,8'h2b,8'h2b,8'h1a,8'h1a,8'h1a,8'h2b,8'h2b,8'h1a,8'h1a,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h1a,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h1a,8'h2b,8'h1a,8'h2b,8'h1a,8'h1a,8'h1a,8'h16,8'h6,8'h6,8'h21,8'h1a,8'h1a,8'h1a,8'h3,8'h6,8'h22,8'h1a,8'h1a,8'h1a,8'h2b,8'h2b,8'h2b,8'h2b,8'h1a,8'h1a,8'h1a,8'h1a,8'h1a,8'h1a,8'h6,8'h6,8'h6,8'h6,8'h6,8'h6,8'h3,8'h1a,8'h1a,8'h1a,8'h1a,8'h1a,8'h1a,8'h2b,8'h1a,8'h1a,8'h2b,8'h1a,8'h1a,8'h1a,8'h0,8'h6,8'h2a,8'h1a,8'h2b,8'h16,8'h22,8'h6,8'h6,8'h1a,8'h1a,8'h1a,8'h1a,8'h1a,8'h1a,8'h1a,8'h1a,8'h1a,8'h1a,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h1a,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h1a,8'h1a,8'h2b,8'h2b,8'h2b,8'h2b,8'h1a,8'h1a,8'h1a,8'h1a,8'h1a,8'h1a,8'h2b,8'h2b,8'h1a,8'h1a,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h1a,8'h1a,8'h1a,8'h1a,8'h1a,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h1a,8'h1a,8'h2b,8'h2b,8'h2b,8'h1a,8'h2b,8'h2b,8'h2b,8'h1a,8'h1a,8'h1a,8'h2b,8'h2b,8'h1a,8'h1a,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h1a,8'h1a,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h1a,8'h1a,8'h1a,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h1a,8'h1a,8'h1a,8'h1a,8'h1a,8'h1a,8'h1a,8'h1a,8'h2b,8'h1a,8'h1a,8'h1a,8'h1a,8'h1a,8'h1a,8'h2b,8'h1a,8'h1a,8'h2b,8'h1a,8'h1a,8'h1a,8'h1a,8'h2b,8'h1a,8'h2b,8'h1a,8'h1a,8'h1a,8'h2b,8'h1a,8'h1a,8'h1a,8'h1a,8'h2b,8'h1a,8'h1a,8'h2b,8'h1a,8'h1a,8'h1a,8'h2b,8'h1a,8'h1a,8'h2b,8'h2b,8'h1a,8'h1a,8'h1a,8'h1a,8'h1a,8'h1a,8'h1a,8'h1a,8'h1a,8'h1a,8'h1a,8'h1a,8'h2b,8'h1a,8'h1a,8'h1a,8'h1a,8'h1a,8'h1a,8'h2b,8'h1a,8'h2b,8'h1a,8'h1a,8'h1a,8'h2b,8'h2b,8'h1a,8'h1a,8'h1a,8'h1a,8'h1a,8'h1a,8'h1a,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h1a,8'h2b,8'h2b,8'h21,8'h6,8'h6,8'h1a,8'h1a,8'h1a,8'h1a,8'h21,8'h6,8'h6,8'h1b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h1a,8'h1a,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h1a,8'h1a,8'h1a,8'h1a,8'h21,8'h6,8'h6,8'h6,8'h6,8'h6,8'h6,8'h21,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h1a,8'h2b,8'h2b,8'h2b,8'h1a,8'h1a,8'h1a,8'h1a,8'h1a,8'h1a,8'h1a,8'h1a,8'h1a,8'h1a,8'h1a,8'h1a,8'h2b,8'h2b,8'h1a,8'h1a,8'h1a,8'h2b,8'h1a,8'h1a,8'h1a,8'h1a,8'h1a,8'h1a,8'h2b,8'h2b,8'h1a,8'h1a,8'h1a,8'h1a,8'h1a,8'h1a,8'h1a,8'h1a,8'h1a,8'h1a,8'h1a,8'h1a,8'h1a,8'h1a,8'h1a,8'h1a,8'h1a,8'h1a,8'h1a,8'h1a,8'h1a,8'h2b,8'h1a,8'h2b,8'h1a,8'h2b,8'h1a,8'h1a,8'h1a,8'h1a,8'h2b,8'h2b,8'h1a,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h1a,8'h2b,8'h2b,8'h2b,8'h1a,8'h21,8'h6,8'h6,8'h1a,8'h1a,8'h1a,8'h2b,8'h1b,8'h22,8'h6,8'h3,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h1a,8'h1a,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h1a,8'h1a,8'h1a,8'h1a,8'h1a,8'h1a,8'h1a,8'h1a,8'h2b,8'h1a,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h1a,8'h2b,8'h2b,8'h2b,8'h1a,8'h1a,8'h1a,8'h1a,8'h1a,8'h1a,8'h1a,8'h9,8'h6,8'h6,8'h6,8'h6,8'h6,8'h1a,8'h1a,8'h2b,8'h2b,8'h1a,8'h2b,8'h1a,8'h2b,8'h1a,8'h2b,8'h2b,8'h1a,8'h1a,8'h2b,8'h1a,8'h1a,8'h1a,8'h1a,8'h1a,8'h1a,8'h2b,8'h1a,8'h1a,8'h1a,8'h1a,8'h1a,8'h1a,8'h1a,8'ha,8'h6,8'h2,8'h1a,8'h1a,8'h1a,8'h1a,8'h2b,8'h2b,8'h1a,8'h1a,8'h2b,8'h2b,8'h2b,8'h1a,8'h1a,8'h1a,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h1a,8'h1a,8'h2b,8'h2b,8'h1a,8'h1a,8'h2b,8'h1a,8'h1a,8'h1a,8'h2b,8'h2b,8'h1a,8'h1a,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h1a,8'h1a,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h1a,8'h1a,8'h1a,8'h1a,8'h1a,8'h1a,8'h2b,8'h2b,8'h2b,8'h2b,8'h1a,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h1a,8'h2b,8'h2b,8'h2b,8'h1a,8'h1a,8'h1a,8'h1a,8'h1a,8'h1a,8'h1a,8'h9,8'h6,8'h1b,8'h1a,8'h1a,8'h1a,8'h2b,8'h1a,8'h2b,8'h2b,8'h1a,8'h1a,8'h1a,8'h2b,8'h1a,8'h1a,8'h1a,8'h1a,8'h1a,8'h2b,8'h2b,8'h1a,8'h1a,8'h1a,8'h1a,8'h1a,8'h2b,8'h1a,8'h1a,8'h1a,8'h1a,8'h1a,8'h1a,8'h1a,8'ha,8'h6,8'h3,8'h1a,8'h1a,8'h1a,8'h2b,8'h1a,8'h2b,8'h2b,8'h2b,8'h1a,8'h1a,8'h1a,8'h2b,8'h2b,8'h1a,8'h2b,8'h1a,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h1a,8'h1a,8'h1a,8'h1a,8'h2b,8'h1a,8'h1a,8'h1a,8'h1a,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h1a,8'h1a,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h1a,8'h1a,8'h1a,8'h1a,8'h1a,8'h2b,8'h2b,8'h1a,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h1a,8'h2b,8'h2b,8'h2b,8'h1a,8'h1a,8'h1a,8'h1a,8'h1a,8'h1a,8'h1a,8'h9,8'h6,8'h1b,8'h1a,8'h1a,8'h1a,8'h1b,8'h6,8'h6,8'h1a,8'h16,8'h22,8'h6,8'h1b,8'h1a,8'h6,8'h6,8'h6,8'h6,8'h21,8'h1a,8'h1a,8'h22,8'h6,8'h6,8'h22,8'h3,8'h9,8'h6,8'h1b,8'h1b,8'h6,8'h2a,8'h1a,8'ha,8'h6,8'h6,8'h6,8'h6,8'h21,8'h1b,8'h6,8'h6,8'h6,8'h6,8'h21,8'h1a,8'h1a,8'h2b,8'h2b,8'h1a,8'h2b,8'h1a,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h1a,8'h1a,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h1a,8'h1a,8'h1a,8'h1a,8'h2b,8'h2b,8'h2b,8'h2b,8'h1a,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h1a,8'h1a,8'h1a,8'h1a,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h1a,8'h2b,8'h2b,8'h2b,8'h1a,8'h1a,8'h2b,8'h2b,8'h1a,8'h1a,8'h1a,8'h9,8'h6,8'h6,8'h6,8'h6,8'h9,8'h1a,8'h1b,8'h6,8'h6,8'h6,8'h6,8'h1a,8'h2b,8'h22,8'h6,8'h1a,8'h2b,8'h6,8'h6,8'h1a,8'h6,8'h6,8'h21,8'h1a,8'h1a,8'h1a,8'h7,8'h6,8'h1b,8'h1b,8'h6,8'h2a,8'h1a,8'ha,8'h6,8'h2,8'h1a,8'h1a,8'h1a,8'h6,8'h22,8'h1a,8'h2b,8'h22,8'h6,8'h1a,8'h2b,8'h1a,8'h1a,8'h1a,8'h2b,8'h1a,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h1a,8'h1a,8'h1a,8'h1a,8'h2b,8'h2b,8'h1a,8'h1a,8'h1a,8'h1a,8'h1a,8'h1a,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h1a,8'h1a,8'h1a,8'h1a,8'h2b,8'h1a,8'h1a,8'h2b,8'h1a,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h1a,8'h2b,8'h2b,8'h2b,8'h1a,8'h1a,8'h2b,8'h2b,8'h1a,8'h1a,8'h1a,8'h9,8'h6,8'h21,8'h1a,8'h1a,8'h2b,8'h2b,8'h1a,8'h21,8'h6,8'h6,8'h1b,8'h2b,8'h1b,8'h6,8'h6,8'h6,8'h6,8'h6,8'h6,8'h3,8'h6,8'h9,8'h1a,8'h1a,8'h1a,8'h1a,8'h6,8'h6,8'h1b,8'h1b,8'h6,8'h2a,8'h1a,8'ha,8'h6,8'h21,8'h1a,8'h1a,8'h1b,8'h6,8'h6,8'h6,8'h6,8'h6,8'h6,8'h1b,8'h2b,8'h1a,8'h2b,8'h2b,8'h2b,8'h1a,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h1a,8'h2b,8'h1a,8'h2b,8'h1a,8'h1a,8'h1a,8'h1a,8'h1a,8'h1a,8'h1a,8'h2b,8'h2b,8'h2b,8'h1a,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h1a,8'h1a,8'h1a,8'h1a,8'h2b,8'h2b,8'h2b,8'h2b,8'h1a,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h1a,8'h2b,8'h2b,8'h2b,8'h1a,8'h1a,8'h2b,8'h2b,8'h1a,8'h1a,8'h1a,8'h9,8'h6,8'h1a,8'h1a,8'h1a,8'h1a,8'h2b,8'h1a,8'h9,8'h6,8'h6,8'h3,8'h2b,8'h1b,8'h6,8'h22,8'h1a,8'h2b,8'h1a,8'h1a,8'h1b,8'h6,8'h22,8'h1a,8'h1a,8'h1a,8'h1a,8'h6,8'h6,8'h1b,8'h1b,8'h6,8'h2a,8'h18,8'h4,8'h6,8'h2,8'h1a,8'h1a,8'h1b,8'h6,8'h22,8'h1a,8'h2b,8'h2b,8'h1a,8'h2b,8'h2b,8'h1a,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h1a,8'h2b,8'h1a,8'h1a,8'h1a,8'h1a,8'h1a,8'h1a,8'h1a,8'h1a,8'h1a,8'h1a,8'h2b,8'h1a,8'h1a,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h1a,8'h1a,8'h1a,8'h1a,8'h2b,8'h1a,8'h1a,8'h2b,8'h2b,8'h1a,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h1a,8'h1a,8'h2b,8'h2b,8'h1a,8'h1a,8'h2b,8'h2b,8'h1a,8'h1a,8'h1a,8'h9,8'h6,8'h1b,8'h1a,8'h1a,8'h2b,8'h2b,8'h3,8'h6,8'h3,8'h2,8'h6,8'h21,8'h1a,8'h6,8'h6,8'h21,8'h1a,8'h2b,8'h1a,8'h1a,8'h6,8'h6,8'h1b,8'h2b,8'h1a,8'h1a,8'h9,8'h6,8'h21,8'h1b,8'h6,8'h2,8'h1a,8'h4,8'h6,8'h2a,8'h1a,8'h1a,8'h1a,8'h22,8'h6,8'h21,8'h2b,8'h1a,8'h2b,8'h1a,8'h2b,8'h2b,8'h1a,8'h2b,8'h2b,8'h1a,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h1a,8'h2b,8'h1a,8'h2b,8'h1a,8'h1a,8'h1a,8'h1a,8'h1a,8'h1a,8'h1a,8'h1a,8'h2b,8'h2b,8'h2b,8'h1a,8'h2b,8'h1a,8'h2b,8'h2b,8'h1a,8'h2b,8'h2b,8'h1a,8'h1a,8'h1a,8'h2b,8'h1a,8'h2b,8'h1a,8'h2b,8'h2b,8'h1a,8'h2b,8'h2b,8'h1a,8'h2b,8'h1a,8'h1a,8'h2b,8'h1a,8'h2b,8'h1a,8'h2b,8'h1a,8'h1a,8'h2b,8'h1a,8'h1a,8'h1a,8'h1a,8'h1a,8'h1a,8'h1a,8'h1a,8'h2b,8'h2b,8'h1a,8'h2b,8'h2b,8'h1a,8'h2b,8'h2b,8'h1a,8'h2b,8'h2b,8'h1a,8'h2b,8'h2b,8'h2b,8'h1a,8'h1a,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h1a,8'h1a,8'h2b,8'h2b,8'h1a,8'h1a,8'h2b,8'h2b,8'h1a,8'h1a,8'h16,8'h3,8'h6,8'h6,8'h6,8'h6,8'h6,8'h6,8'h6,8'h9,8'h1a,8'h1b,8'h6,8'h6,8'h21,8'h1b,8'h6,8'h6,8'h6,8'h6,8'h2,8'h1a,8'h1a,8'h6,8'h6,8'h6,8'h6,8'h21,8'h16,8'h6,8'h6,8'h6,8'h6,8'h2,8'h1a,8'h1a,8'h2,8'h6,8'h6,8'h6,8'h3,8'h16,8'h6,8'h6,8'h6,8'h6,8'h2,8'h1a,8'h2b,8'h1a,8'h1a,8'h2b,8'h1a,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h1a,8'h1a,8'h1a,8'h2b,8'h1a,8'h1a,8'h1a,8'h1a,8'h1a,8'h1a,8'h1a,8'h1a,8'h2b,8'h1a,8'h1a,8'h2b,8'h1a,8'h2b,8'h2b,8'h1a,8'h2b,8'h1a,8'h1a,8'h2b,8'h1a,8'h1a,8'h1a,8'h1a,8'h2b,8'h2b,8'h1a,8'h2b,8'h2b,8'h1a,8'h1a,8'h2b,8'h2b,8'h1a,8'h2b,8'h2b,8'h1a,8'h1a,8'h1a,8'h2b,8'h2b,8'h2b,8'h1a,8'h2b,8'h16,8'h1a,8'h1a,8'h2b,8'h1a,8'h2b,8'h2b,8'h1a,8'h1a,8'h2b,8'h2b,8'h1a,8'h2b,8'h2b,8'h2b,8'h2b,8'h1a,8'h1a,8'h1a,8'h2b,8'h2b,8'h1a,8'h1a,8'h2b,8'h2b,8'h1a,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h1a,8'h1a,8'h2b,8'h2b,8'h1a,8'h1a,8'h2b,8'h2b,8'h1a,8'h1a,8'h1a,8'h1a,8'h1a,8'h1a,8'h2b,8'h1a,8'h1a,8'h1a,8'h2b,8'h2b,8'h2b,8'h1a,8'h1a,8'h1a,8'h1a,8'h2b,8'h1a,8'h2b,8'h1a,8'h1a,8'h2b,8'h2b,8'h1a,8'h2b,8'h2b,8'h1a,8'h1a,8'h2b,8'h1a,8'h1a,8'h1a,8'h1a,8'h1a,8'h1a,8'h1a,8'h1a,8'h1a,8'h1a,8'h1a,8'h1a,8'h1a,8'h2b,8'h1a,8'h1a,8'h1a,8'h2b,8'h1a,8'h2b,8'h1a,8'h1a,8'h2b,8'h2b,8'h1a,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h1a,8'h1a,8'h1a,8'h1a,8'h1a,8'h1a,8'h1a,8'h1a,8'h1a,8'h1a,8'h1a,8'h1a,8'h2b,8'h1a,8'h2b,8'h2b,8'h1a,8'h2b,8'h1a,8'h1a,8'h2b,8'h2b,8'h2b,8'h1a,8'h1a,8'h1a,8'h2b,8'h2b,8'h1a,8'h1a,8'h1a,8'h1a,8'h1a,8'h2b,8'h2b,8'h1a,8'h1a,8'h2b,8'h1a,8'h1a,8'h1a,8'h2b,8'h1a,8'h2b,8'h1a,8'h1a,8'h2b,8'h1a,8'h2b,8'h1a,8'h1a,8'h2b,8'h2b,8'h2b,8'h1a,8'h2b,8'h2b,8'h1a,8'h1a,8'h2b,8'h1a,8'h1a,8'h1a,8'h1a,8'h2b,8'h2b,8'h2b,8'h2b,8'h1a,8'h1a,8'h1a,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h1a,8'h1a,8'h2b,8'h2b,8'h1a,8'h1a,8'h2b,8'h2b,8'h2b,8'h1a,8'h1a,8'h1a,8'h2b,8'h2b,8'h1a,8'h1a,8'h1a,8'h1a,8'h2b,8'h2b,8'h1a,8'h1a,8'h1a,8'h1a,8'h2b,8'h1a,8'h1a,8'h2b,8'h1a,8'h1a,8'h2b,8'h1a,8'h2b,8'h2b,8'h1a,8'h1a,8'h1a,8'h1a,8'h1a,8'h1a,8'h2b,8'h2b,8'h1a,8'h1a,8'h1a,8'h1a,8'h1a,8'h1a,8'h1a,8'h1a,8'h1a,8'h1a,8'h2b,8'h2b,8'h1a,8'h2b,8'h2b,8'h2b,8'h1a,8'h1a,8'h2b,8'h2b,8'h1a,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h1a,8'h1a,8'h1a,8'h1a,8'h1a,8'h1a,8'h1a,8'h1a,8'ha,8'h6,8'h21,8'h2b,8'h1a,8'h2b,8'h3,8'h6,8'h1b,8'h1a,8'h2b,8'h1a,8'h1a,8'h1a,8'h2b,8'h2b,8'h1a,8'h1a,8'h1a,8'h1a,8'h2b,8'h2b,8'h2b,8'h2b,8'h1a,8'h2b,8'h1a,8'h1a,8'h1a,8'h2b,8'h2b,8'h2b,8'h1a,8'h2b,8'h2b,8'h1a,8'h1a,8'h2b,8'h2b,8'h1a,8'h1a,8'h2b,8'h2b,8'h1a,8'h2b,8'h2b,8'h2b,8'h2b,8'h1a,8'h2b,8'h2b,8'h2b,8'h1a,8'h2b,8'h21,8'h6,8'h21,8'h1a,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h1a,8'h1a,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h1a,8'h1a,8'h2b,8'h2b,8'h1a,8'h1a,8'h2b,8'h2b,8'h1a,8'h1a,8'h1a,8'h1a,8'h1a,8'h2b,8'h2b,8'h1a,8'h1a,8'h1a,8'h1a,8'h2b,8'h2b,8'h2b,8'h1a,8'h1a,8'h2b,8'h2b,8'h2b,8'h1a,8'h2b,8'h1a,8'h2b,8'h2b,8'h1a,8'h1a,8'h1a,8'h2b,8'h1a,8'h1a,8'h1a,8'h1a,8'h1a,8'h1a,8'h1a,8'h1a,8'h1a,8'h1a,8'h2b,8'h1a,8'h1a,8'h1a,8'h1a,8'h1a,8'h1a,8'h1a,8'h2b,8'h1a,8'h1a,8'h1a,8'h2b,8'h2b,8'h1a,8'h1a,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h1a,8'h1a,8'h1a,8'h1a,8'h1a,8'h1a,8'h1a,8'h1a,8'h3,8'h6,8'h3,8'h1a,8'h1a,8'h16,8'h6,8'h6,8'h21,8'h1a,8'h1a,8'h2b,8'h1a,8'h2b,8'h1a,8'h2b,8'h1a,8'h1a,8'h1a,8'h1a,8'h1a,8'h1a,8'h2b,8'h2b,8'h1a,8'h2b,8'h1a,8'h2b,8'h2b,8'h1a,8'h1a,8'h2b,8'h1a,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h1a,8'h1a,8'h1a,8'h1a,8'h1a,8'h2b,8'h2b,8'h1a,8'h1a,8'h2b,8'h1a,8'h2b,8'h1a,8'h2b,8'h1a,8'h3,8'h6,8'h21,8'h1a,8'h1a,8'h1a,8'h1a,8'h1a,8'h2b,8'h2b,8'h2b,8'h1a,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h1a,8'h1a,8'h2b,8'h2b,8'h1a,8'h1a,8'h2b,8'h2b,8'h1a,8'h1a,8'h1a,8'h1a,8'h1a,8'h1a,8'h2b,8'h1a,8'h2b,8'h2b,8'h1a,8'h1a,8'h2b,8'h1a,8'h1a,8'h2b,8'h1a,8'h1a,8'h1a,8'h1a,8'h2b,8'h2b,8'h1a,8'h1a,8'h1a,8'h2b,8'h1a,8'h1a,8'h1a,8'h1a,8'h1a,8'h1a,8'h1a,8'h2b,8'h1a,8'h1a,8'h1a,8'h1a,8'h2b,8'h1a,8'h1a,8'h1a,8'h1a,8'h2b,8'h1a,8'h1a,8'h2b,8'h2b,8'h1a,8'h2b,8'h2b,8'h1a,8'h1a,8'h2b,8'h2b,8'h1a,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h1a,8'h1a,8'h1a,8'h1a,8'h1a,8'h1a,8'h1a,8'h1a,8'h9,8'h6,8'h6,8'h1b,8'h2b,8'h3,8'h6,8'h6,8'h21,8'h1a,8'h1b,8'h6,8'h6,8'h6,8'h6,8'h1b,8'h21,8'h6,8'h21,8'h1a,8'h3,8'h6,8'h1b,8'h1b,8'h22,8'h6,8'h6,8'h6,8'h21,8'h1a,8'h9,8'h6,8'h6,8'h6,8'h6,8'h6,8'h6,8'h6,8'h21,8'h1a,8'h1a,8'h22,8'h6,8'h6,8'h6,8'h21,8'h1a,8'h22,8'h6,8'h6,8'h6,8'h6,8'h1a,8'h2b,8'h3,8'h6,8'h6,8'h6,8'h6,8'h21,8'h2b,8'h2b,8'h1a,8'h1a,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h1a,8'h1a,8'h2b,8'h2b,8'h1a,8'h1a,8'h2b,8'h2b,8'h2b,8'h1a,8'h1a,8'h1a,8'h2b,8'h2b,8'h2b,8'h1a,8'h1a,8'h1a,8'h1a,8'h1a,8'h2b,8'h2b,8'h2b,8'h1a,8'h1a,8'h1a,8'h1a,8'h1a,8'h2b,8'h2b,8'h2b,8'h1a,8'h1a,8'h2b,8'h1a,8'h1a,8'h2b,8'h1a,8'h2b,8'h1a,8'h1a,8'h1a,8'h1a,8'h1a,8'h1a,8'h1a,8'h2b,8'h1a,8'h1a,8'h1a,8'h1a,8'h2b,8'h2b,8'h2b,8'h1a,8'h2b,8'h2b,8'h1a,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h1a,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h1a,8'h1a,8'h1a,8'h1a,8'h1a,8'h1a,8'h1a,8'h1a,8'h9,8'h9,8'h3,8'h3,8'h16,8'h6,8'h6,8'h6,8'h3,8'h1a,8'h22,8'h6,8'h1b,8'h16,8'h6,8'h9,8'h21,8'h6,8'h9,8'h1a,8'h6,8'h22,8'h1b,8'h22,8'h6,8'h16,8'h1a,8'h22,8'h6,8'h16,8'h6,8'h6,8'h16,8'h9,8'h6,8'h21,8'h1a,8'h9,8'h9,8'h1a,8'h22,8'h6,8'h1a,8'h2b,8'h6,8'h6,8'h1a,8'h22,8'h6,8'h1b,8'h1b,8'h6,8'h2,8'h1a,8'h3,8'h6,8'h3,8'h2b,8'h1a,8'h2b,8'h2b,8'h1a,8'h1a,8'h2b,8'h2b,8'h1a,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h1a,8'h1a,8'h2b,8'h2b,8'h1a,8'h1a,8'h2b,8'h2b,8'h2b,8'h1a,8'h1a,8'h1a,8'h2b,8'h2b,8'h2b,8'h1a,8'h1a,8'h2b,8'h2b,8'h2b,8'h1a,8'h1a,8'h2b,8'h2b,8'h2b,8'h1a,8'h1a,8'h2b,8'h2b,8'h2b,8'h2b,8'h1a,8'h1a,8'h1a,8'h1a,8'h1a,8'h1a,8'h1a,8'h2b,8'h1a,8'h1a,8'h1a,8'h1a,8'h1a,8'h1a,8'h1a,8'h1a,8'h1a,8'h1a,8'h1a,8'h1a,8'h1a,8'h2b,8'h1a,8'h1a,8'h2b,8'h1a,8'h1a,8'h2b,8'h2b,8'h2b,8'h1a,8'h1a,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h1a,8'h1a,8'h1a,8'h1a,8'h1a,8'h1a,8'h1a,8'h16,8'h6,8'h9,8'h21,8'h6,8'h6,8'h6,8'h6,8'h6,8'h9,8'h1b,8'h6,8'h2,8'h2b,8'h1a,8'h6,8'h6,8'h1b,8'h22,8'h6,8'h21,8'h6,8'h2,8'h1b,8'h6,8'h6,8'h6,8'h6,8'h6,8'h6,8'h1b,8'h6,8'h6,8'h2b,8'h21,8'h6,8'h3,8'h2b,8'h21,8'h3,8'h1b,8'h6,8'h6,8'h6,8'h6,8'h6,8'h6,8'h1b,8'h22,8'h6,8'h1b,8'h1a,8'h2,8'h3,8'h2b,8'h3,8'h6,8'h21,8'h1a,8'h2b,8'h2b,8'h1a,8'h2b,8'h2b,8'h1a,8'h1a,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h1a,8'h1a,8'h2b,8'h2b,8'h1a,8'h1a,8'h2b,8'h2b,8'h1a,8'h1a,8'h1a,8'h1a,8'h2b,8'h2b,8'h2b,8'h1a,8'h1a,8'h2b,8'h1a,8'h1a,8'h2b,8'h1a,8'h1a,8'h1a,8'h2b,8'h2b,8'h1a,8'h2b,8'h1a,8'h1a,8'h2b,8'h2b,8'h1a,8'h2b,8'h1a,8'h1a,8'h1a,8'h1a,8'h2b,8'h2b,8'h1a,8'h1a,8'h1a,8'h1a,8'h1a,8'h1a,8'h2b,8'h1a,8'h1a,8'h1a,8'h1a,8'h1a,8'h2b,8'h2b,8'h2b,8'h1a,8'h2b,8'h2b,8'h1a,8'h1a,8'h1a,8'h2b,8'h1a,8'h1a,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h1a,8'h2b,8'h1a,8'h2b,8'h1a,8'h6,8'h22,8'h1b,8'h22,8'h6,8'h9,8'h16,8'h6,8'h9,8'h1b,8'h6,8'h2,8'h1a,8'h1a,8'h22,8'h6,8'h1b,8'h3,8'h6,8'h6,8'h6,8'h1b,8'h1b,8'h6,8'h22,8'h1a,8'h2b,8'h1a,8'h1a,8'h1a,8'h6,8'h6,8'h1a,8'h21,8'h6,8'h3,8'h2b,8'h3,8'h3,8'h1b,8'h6,8'h22,8'h1a,8'h1a,8'h1a,8'h1a,8'h1a,8'h6,8'h6,8'h1b,8'h1a,8'h9,8'h9,8'h16,8'h21,8'h6,8'h3,8'h1a,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h1a,8'h1a,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h1a,8'h2b,8'h2b,8'h1a,8'h1a,8'h2b,8'h1a,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h1a,8'h1a,8'h2b,8'h2b,8'h2b,8'h1a,8'h1a,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h1a,8'h2b,8'h2b,8'h1a,8'h1a,8'h2b,8'h2b,8'h1a,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h1a,8'h2b,8'h2b,8'h2b,8'h1a,8'h1a,8'h2b,8'h2b,8'h1a,8'h2b,8'h2b,8'h2b,8'h1a,8'h1a,8'h2b,8'h2b,8'h1a,8'h1a,8'h1a,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h1a,8'h2b,8'h2b,8'h1a,8'h2b,8'h1a,8'h1a,8'h2b,8'h2b,8'h2b,8'h1a,8'h2b,8'h2b,8'h2b,8'h1a,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h1a,8'h1a,8'h1b,8'h6,8'h9,8'h1a,8'h9,8'h6,8'h21,8'h1a,8'h6,8'h9,8'h1a,8'h22,8'h6,8'h1b,8'h1b,8'h6,8'h9,8'h1a,8'h1b,8'h6,8'h6,8'h9,8'h2b,8'h1a,8'h6,8'h6,8'h21,8'h2b,8'h2b,8'h1a,8'h1a,8'h22,8'h6,8'h1a,8'h21,8'h6,8'h3,8'h2b,8'h21,8'h3,8'h1b,8'h22,8'h6,8'h21,8'h1a,8'h2b,8'h1a,8'h2b,8'h22,8'h6,8'h1b,8'h1a,8'h9,8'h9,8'h1a,8'h21,8'h6,8'h9,8'h2b,8'h1a,8'h1a,8'h2b,8'h1a,8'h2b,8'h2b,8'h2b,8'h1a,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h1a,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h1a,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h1a,8'h1a,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h1a,8'h1a,8'h2b,8'h2b,8'h2b,8'h1a,8'h1a,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h1a,8'h1a,8'h2b,8'h2b,8'h2b,8'h2b,8'h1a,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h1a,8'h1a,8'h1a,8'h2b,8'h2b,8'h2b,8'h2b,8'h1a,8'h1a,8'h1a,8'h2b,8'h2b,8'h2b,8'h2b,8'h1a,8'h1a,8'h1a,8'h1a,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h1a,8'h1a,8'h1a,8'h1a,8'h1a,8'h1a,8'h1a,8'h1a,8'h1a,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h1a,8'h1a,8'h2b,8'h2b,8'h1a,8'h1b,8'h22,8'h22,8'h1a,8'h1a,8'h1a,8'h2b,8'h1b,8'h6,8'h9,8'h1a,8'h1a,8'h6,8'h6,8'h6,8'h6,8'h1a,8'h2b,8'h1a,8'h2,8'h6,8'h21,8'h1a,8'h1a,8'h16,8'h6,8'h6,8'h6,8'h6,8'h3,8'h1a,8'h6,8'h6,8'h1a,8'h21,8'h6,8'h21,8'h1a,8'h3,8'h2,8'h1a,8'h1b,8'h6,8'h6,8'h6,8'h6,8'h2,8'h1a,8'h22,8'h6,8'h1b,8'h1a,8'h9,8'h9,8'h1a,8'h1a,8'h9,8'h6,8'h6,8'h6,8'h21,8'h1a,8'h2b,8'h1a,8'h1a,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h1a,8'h1a,8'h1a,8'h1a,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h1a,8'h1a,8'h1a,8'h1a,8'h1a,8'h2b,8'h1a,8'h1a,8'h2b,8'h2b,8'h2b,8'h1a,8'h2b,8'h1a,8'h1a,8'h1a,8'h1a,8'h2b,8'h2b,8'h2b,8'h1a,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h1a,8'h1a,8'h2b,8'h2b,8'h2b,8'h1a,8'h1a,8'h1a,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h1a,8'h1a,8'h2b,8'h2b,8'h1a,8'h1a,8'h2b,8'h2b,8'h1a,8'h1a,8'h2b,8'h2b,8'h2b,8'h2b,8'h1a,8'h1a,8'h1a,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h1a,8'h1a,8'h2b,8'h2b,8'h2b,8'h1a,8'h1a,8'h1a,8'h2b,8'h2b,8'h2b,8'h2b,8'h1a,8'h1a,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h1a,8'h1a,8'h1a,8'h2b,8'h1a,8'h2b,8'h1a,8'h2b,8'h1a,8'h1a,8'h1a,8'h1a,8'h1a,8'h2b,8'h2b,8'h2b,8'h1a,8'h1a,8'h1a,8'h2b,8'h1a,8'h1a,8'h1a,8'h2b,8'h1a,8'h2b,8'h1a,8'h1a,8'h2b,8'h1a,8'h2b,8'h2b,8'h1a,8'h1a,8'h2b,8'h1a,8'h1a,8'h1a,8'h1a,8'h1a,8'h2b,8'h1a,8'h2b,8'h2b,8'h2b,8'h1a,8'h1a,8'h1a,8'h1a,8'h1a,8'h2b,8'h2b,8'h2b,8'h2b,8'h1a,8'h1a,8'h1a,8'h2b,8'h2b,8'h1a,8'h2b,8'h1a,8'h1a,8'h1a,8'h1a,8'h1a,8'h2b,8'h2b,8'h2b,8'h1a,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h1a,8'h1a,8'h2b,8'h2b,8'h1a,8'h1a,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h1a,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h1a,8'h1a,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h1a,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h1a,8'h1a,8'h2b,8'h2b,8'h1a,8'h1a,8'h1a,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h1a,8'h1a,8'h2b,8'h1a,8'h2b,8'h1a,8'h1a,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h1a,8'h1a,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h1a,8'h2b,8'h2b,8'h1a,8'h1a,8'h2b,8'h1a,8'h2b,8'h2b,8'h1a,8'h1a,8'h1a,8'h2b,8'h2b,8'h1a,8'h2b,8'h1a,8'h1a,8'h2b,8'h1a,8'h2b,8'h1a,8'h1a,8'h1a,8'h1a,8'h1a,8'h1a,8'h1a,8'h2b,8'h1a,8'h1a,8'h1a,8'h1a,8'h1a,8'h2b,8'h2b,8'h1a,8'h1a,8'h2b,8'h2b,8'h1a,8'h1a,8'h2b,8'h1a,8'h2b,8'h1a,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h1a,8'h1a,8'h2b,8'h1a,8'h1a,8'h1a,8'h1a,8'h1a,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h1a,8'h1a,8'h1a,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h1a,8'h1a,8'h2b,8'h2b,8'h2b,8'h2b,8'h1a,8'h1a,8'h1a,8'h2b,8'h2b,8'h1a,8'h1a,8'h1a,8'h2b,8'h2b,8'h2b,8'h2b,8'h1a,8'h2b,8'h1a,8'h1a,8'h1a,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h1a,8'h1a,8'h2b,8'h2b,8'h2b,8'h1a,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h1a,8'h1a,8'h1a,8'h1a,8'h1a,8'h1a,8'h1a,8'h1a,8'h1a,8'h1a,8'h2b,8'h2b,8'h2b,8'h2b,8'h1a,8'h2b,8'h1a,8'h1a,8'h1a,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h1a,8'h1a,8'h2b,8'h1a,8'h1a,8'h1a,8'h1a,8'h2b,8'h1a,8'h1a,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h1a,8'h2b,8'h1a,8'h1a,8'h2b,8'h2b,8'h1a,8'h1a,8'h1a,8'h1a,8'h1a,8'h1a,8'h1a,8'h1a,8'h2b,8'h1a,8'h1a,8'h1a,8'h1a,8'h2b,8'h2b,8'h1a,8'h1a,8'h1a,8'h2b,8'h2b,8'h1a,8'h1a,8'h1a,8'h2b,8'h2b,8'h2b,8'h1a,8'h1a,8'h2b,8'h2b,8'h1a,8'h1a,8'h1a,8'h2b,8'h1a,8'h2b,8'h2b,8'h1a,8'h1a,8'h2b,8'h2b,8'h1a,8'h2b,8'h2b,8'h1a,8'h2b,8'h2b,8'h1a,8'h1a,8'h1a,8'h2b,8'h2b,8'h2b,8'h1a,8'h1a,8'h1a,8'h2b,8'h1a,8'h1a,8'h1a,8'h2b,8'h1a,8'h1a,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h1a,8'h2b,8'h2b,8'h1a,8'h1a,8'h2b,8'h2b,8'h1a,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h1a,8'h1a,8'h2b,8'h2b,8'h1a,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h1a,8'h1a,8'h2b,8'h2b,8'h2b,8'h1a,8'h1a,8'h1a,8'h2b,8'h2b,8'h2b,8'h1a,8'h1a,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h1a,8'h2b,8'h2b,8'h2b,8'h1a,8'h1a,8'h1a,8'h1a,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h1a,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h1a,8'h2b,8'h2b,8'h2b,8'h1a,8'h1a,8'h1a,8'h1a,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h1a,8'h2b,8'h2b,8'h2b,8'h1a,8'h1a,8'h1a,8'h2b,8'h2b,8'h2b,8'h2b,8'h1a,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h1a,8'h2b,8'h2b,8'h1a,8'h1a,8'h1a,8'h1a,8'h1a,8'h1a,8'h1a,8'h2b,8'h2b,8'h2b,8'h1a,8'h2b,8'h2b,8'h1a,8'h2b,8'h1a,8'h1a,8'h2b,8'h2b,8'h1a,8'h1a,8'h1a,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h1a,8'h1a,8'h2b,8'h1a,8'h2b,8'h1a,8'h1a,8'h2b,8'h1a,8'h2b,8'h2b,8'h2b,8'h2b,8'h1a,8'h2b,8'h1a,8'h2b,8'h1a,8'h2b,8'h2b,8'h1a,8'h2b,8'h1a,8'h1a,8'h2b,8'h1a,8'h1a,8'h1a,8'h1a,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h1a,8'h2b,8'h2b,8'h1a,8'h1a,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h1a,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h1a,8'h1a,8'h2b,8'h2b,8'h1a,8'h1a,8'h2b,8'h2b,8'h1a,8'h1a,8'h2b,8'h2b,8'h2b,8'h1a,8'h1a,8'h1a,8'h2b,8'h2b,8'h1a,8'h1a,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h1a,8'h1a,8'h2b,8'h2b,8'h1a,8'h1a,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h1a,8'h2b,8'h2b,8'h2b,8'h1a,8'h1a,8'h1a,8'h2b,8'h1a,8'h1a,8'h2b,8'h1a,8'h1a,8'h2b,8'h2b,8'h2b,8'h1a,8'h1a,8'h1a,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h1a,8'h1a,8'h1a,8'h1a,8'h1a,8'h1a,8'h1a,8'h1a,8'h2b,8'h2b,8'h2b,8'h1a,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h1a,8'h2b,8'h2b,8'h2b,8'h2b,8'h1a,8'h2b,8'h2b,8'h2b,8'h1a,8'h2b,8'h1a,8'h2b,8'h2b,8'h2b,8'h1a,8'h2b,8'h2b,8'h1a,8'h2b,8'h2b,8'h1a,8'h2b,8'h1a,8'h1a,8'h2b,8'h2b,8'h2b,8'h1a,8'h2b,8'h1a,8'h2b,8'h2b,8'h2b,8'h2b,8'h1a,8'h2b,8'h2b,8'h1a,8'h2b,8'h2b,8'h1a,8'h2b,8'h1a,8'h2b,8'h2b,8'h1a,8'h1a,8'h2b,8'h1a,8'h2b,8'h2b,8'h1a,8'h2b,8'h2b,8'h2b,8'h2b,8'h1a,8'h1a,8'h1a,8'h2b,8'h1a,8'h2b,8'h2b,8'h2b,8'h1a,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h1a,8'h21,8'h3,8'h21,8'h3,8'h3,8'h21,8'h1a,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h1a,8'h2b,8'h2b,8'h1a,8'h21,8'h21,8'h3,8'h21,8'h3,8'h21,8'h16,8'h2b,8'h2b,8'h1a,8'h2b,8'h1a,8'h2b,8'h1a,8'h21,8'h21,8'h1b,8'h1a,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h21,8'h21,8'h1b,8'h1a,8'h2b,8'h1a,8'h1a,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h1a,8'h2b,8'h2b,8'h16,8'h21,8'h3,8'h3,8'h21,8'h21,8'h1b,8'h2b,8'h2b,8'h1a,8'h2b,8'h2b,8'h2b,8'h1a,8'h1a,8'h1a,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h21,8'h21,8'h1b,8'h1a,8'h2b,8'h1a,8'h1b,8'h3,8'h1b,8'h1a,8'h2b,8'h2b,8'h1a,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h21,8'h21,8'h1b,8'h2b,8'h16,8'h3,8'h21,8'h1a,8'h2b,8'h1a,8'h1a,8'h2b,8'h1a,8'h2b,8'h1a,8'h2b,8'h1a,8'h1a,8'h2b,8'h1a,8'h1a,8'h2b,8'h2b,8'h1a,8'h2b,8'h2b,8'h1a,8'h2b,8'h2b,8'h1a,8'h2b,8'h2b,8'h2b,8'h1a,8'h1a,8'h2b,8'h21,8'h3,8'h1a,8'h1a,8'h2b,8'h1a,8'h1a,8'h1a,8'h2b,8'h1a,8'h2b,8'h2b,8'h2b,8'h1a,8'h1b,8'h3,8'h1b,8'h2b,8'h1a,8'h2b,8'h2b,8'h2b,8'h2b,8'h1a,8'h1a,8'h1a,8'h1a,8'h2b,8'h1a,8'h2b,8'h1a,8'h2b,8'h2b,8'h2b,8'h1a,8'h1a,8'h21,8'h3,8'h1b,8'h1a,8'h1a,8'h2b,8'h1a,8'h2b,8'h1a,8'h2b,8'h1a,8'h2b,8'h2b,8'h1a,8'h2b,8'h2b,8'h1a,8'h1a,8'h3,8'h3,8'h1a,8'h1a,8'h2b,8'h2b,8'h1a,8'h2b,8'h1a,8'h2b,8'h1a,8'h2b,8'h2b,8'h1a,8'h1a,8'h1a,8'h2b,8'h1a,8'h2b,8'h2b,8'h1a,8'h21,8'h21,8'h1b,8'h2b,8'h2b,8'h1a,8'h1a,8'h1a,8'h2b,8'h2b,8'h1a,8'h2b,8'h2b,8'h1a,8'h2b,8'h1a,8'h1a,8'h2b,8'h2b,8'h2b,8'h1a,8'h1a,8'h2b,8'h1a,8'h1a,8'h2b,8'h2b,8'h1a,8'h1a,8'h1a,8'h2b,8'h1a,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h1a,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h1a,8'h2b,8'h2b,8'h2b,8'h2b,8'h1a,8'h1a,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h1a,8'h21,8'h21,8'h1b,8'h2b,8'h2b,8'h21,8'h21,8'h1a,8'h21,8'h21,8'h21,8'h3,8'h1b,8'h1a,8'h21,8'h3,8'h21,8'h21,8'h1b,8'h2b,8'h1b,8'h3,8'h3,8'h3,8'h21,8'h1a,8'h21,8'h3,8'h3,8'h3,8'h21,8'h2b,8'h2b,8'h1a,8'h1a,8'h1a,8'h21,8'h21,8'h1b,8'h2b,8'h1a,8'h1a,8'h2b,8'h21,8'h3,8'h21,8'h3,8'h21,8'h1a,8'h2b,8'h21,8'h21,8'h3,8'h3,8'h21,8'h1b,8'h16,8'h21,8'h3,8'h21,8'h21,8'h1b,8'h2b,8'h21,8'h3,8'h3,8'h3,8'h21,8'h1a,8'h2b,8'h2b,8'h1a,8'h1b,8'h3,8'h21,8'h4,8'h21,8'h1b,8'h1a,8'h21,8'h3,8'h3,8'h21,8'h1b,8'h2b,8'h1a,8'h1a,8'h2b,8'h1a,8'h21,8'h21,8'h1b,8'h2b,8'h2b,8'h1a,8'h1a,8'h2b,8'h1b,8'h3,8'h21,8'h3,8'h21,8'h1a,8'h1a,8'h21,8'h3,8'h3,8'h3,8'h21,8'h1b,8'h2b,8'h21,8'h21,8'h21,8'h3,8'h21,8'h1b,8'h1b,8'h4,8'h1b,8'h1a,8'h21,8'h3,8'h21,8'h3,8'h21,8'h1a,8'h1a,8'h21,8'h3,8'h16,8'h16,8'h21,8'h21,8'h2b,8'h1a,8'h3,8'h3,8'h3,8'h21,8'h1b,8'h2b,8'h1a,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h1a,8'h1a,8'h2b,8'h2b,8'h2b,8'h2b,8'h1a,8'h2b,8'h2b,8'h2b,8'h1a,8'h1a,8'h2b,8'h2b,8'h2b,8'h2b,8'h1a,8'h1a,8'h2b,8'h2b,8'h2b,8'h2b,8'h1a,8'h2b,8'h2b,8'h2b,8'h1a,8'h1a,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h1a,8'h1a,8'h1a,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h21,8'h21,8'h1b,8'h1a,8'h1a,8'h3,8'h3,8'h1a,8'h21,8'h3,8'h1b,8'h2b,8'h1a,8'h21,8'h3,8'h1a,8'h1a,8'h21,8'h3,8'h16,8'h21,8'h21,8'h2b,8'h2b,8'h1a,8'h2b,8'h21,8'h21,8'h2b,8'h2b,8'h1a,8'h1a,8'h1a,8'h2b,8'h2b,8'h2b,8'h21,8'h3,8'h21,8'h21,8'h3,8'h21,8'h1a,8'h21,8'h21,8'h1a,8'h1a,8'h3,8'h1b,8'h2b,8'h21,8'h21,8'h21,8'h1a,8'h2b,8'h1a,8'h21,8'h21,8'h1a,8'h1a,8'h21,8'h21,8'h1a,8'h21,8'h21,8'h1a,8'h2b,8'h2b,8'h2b,8'h1a,8'h1a,8'h1a,8'h21,8'h3,8'h1b,8'h1a,8'h2b,8'h1a,8'h21,8'h3,8'h16,8'h16,8'h21,8'h21,8'h1a,8'h2b,8'h1a,8'h1a,8'h1a,8'h3,8'h21,8'h1a,8'h1a,8'h1a,8'h2b,8'h2b,8'h2b,8'h21,8'h3,8'h1a,8'h1a,8'h3,8'h21,8'h1a,8'h21,8'h4,8'h16,8'h1a,8'h21,8'h21,8'h2b,8'h1b,8'h3,8'h21,8'h1a,8'h1a,8'h2b,8'h1b,8'h3,8'h1b,8'h1a,8'h21,8'h3,8'h1a,8'h16,8'h3,8'h21,8'h2b,8'h21,8'h3,8'h1a,8'h1a,8'h3,8'h21,8'h2b,8'h21,8'h21,8'h1a,8'h1a,8'h21,8'h3,8'h16,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h1a,8'h1a,8'h2b,8'h2b,8'h2b,8'h1a,8'h1a,8'h2b,8'h2b,8'h2b,8'h1a,8'h1a,8'h2b,8'h2b,8'h2b,8'h1a,8'h1a,8'h1a,8'h2b,8'h2b,8'h2b,8'h1a,8'h1a,8'h2b,8'h2b,8'h2b,8'h1a,8'h1a,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h1a,8'h1a,8'h1a,8'h1a,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h1a,8'h21,8'h3,8'h21,8'h3,8'h3,8'h21,8'h1a,8'h1a,8'h21,8'h3,8'h1a,8'h2b,8'h1a,8'h3,8'h21,8'h21,8'h3,8'h21,8'h21,8'h1b,8'h21,8'h21,8'h21,8'h1a,8'h2b,8'h1a,8'h21,8'h21,8'h21,8'h1a,8'h2b,8'h2b,8'h2b,8'h1a,8'h1a,8'h1a,8'h21,8'h21,8'h16,8'h1a,8'h2b,8'h1a,8'h2b,8'h21,8'h21,8'h1a,8'h1a,8'h21,8'h21,8'h2b,8'h21,8'h21,8'h1b,8'h2b,8'h1a,8'h1b,8'h21,8'h21,8'h3,8'h3,8'h21,8'h21,8'h16,8'h21,8'h3,8'h1a,8'h1a,8'h1a,8'h1a,8'h1a,8'h2b,8'h1a,8'h21,8'h21,8'h1b,8'h1a,8'h1a,8'h1a,8'h3,8'h21,8'h2b,8'h1a,8'h21,8'h21,8'h1a,8'h1a,8'h2b,8'h1a,8'h1a,8'h3,8'h21,8'h1a,8'h2b,8'h2b,8'h1a,8'h1a,8'h1b,8'h21,8'h21,8'h1a,8'h1a,8'h21,8'h21,8'h1a,8'h21,8'h3,8'h1a,8'h1a,8'h21,8'h21,8'h2b,8'h21,8'h3,8'h1b,8'h2b,8'h1a,8'h1a,8'h1b,8'h3,8'h1b,8'h2b,8'h21,8'h3,8'h16,8'h1a,8'h21,8'h21,8'h1a,8'h21,8'h21,8'h16,8'h1b,8'h21,8'h21,8'h1a,8'h3,8'h3,8'h21,8'h3,8'h3,8'h21,8'h1a,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h1a,8'h1a,8'h2b,8'h2b,8'h2b,8'h1a,8'h1a,8'h2b,8'h2b,8'h2b,8'h1a,8'h1a,8'h2b,8'h2b,8'h2b,8'h1a,8'h1a,8'h1a,8'h2b,8'h2b,8'h2b,8'h1a,8'h1a,8'h2b,8'h2b,8'h2b,8'h1a,8'h1a,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h1a,8'h1a,8'h1a,8'h1a,8'h1a,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h21,8'h3,8'h1b,8'h1a,8'h2b,8'h1a,8'h1a,8'h1a,8'h1b,8'h21,8'h1b,8'h1a,8'h16,8'h3,8'h21,8'h1a,8'h2b,8'h2b,8'h1a,8'h2b,8'h2b,8'h1a,8'h21,8'h3,8'h21,8'h1a,8'h2b,8'h1a,8'h3,8'h3,8'h21,8'h1a,8'h2b,8'h2b,8'h1a,8'h2b,8'h21,8'h3,8'h16,8'h2b,8'h2b,8'h1a,8'h1a,8'h21,8'h3,8'h1a,8'h1a,8'h21,8'h21,8'h1a,8'h21,8'h21,8'h21,8'h1a,8'h2b,8'h1a,8'h3,8'h21,8'h1a,8'h1a,8'h2b,8'h1a,8'h2b,8'h21,8'h3,8'h1a,8'h1a,8'h2b,8'h2b,8'h1a,8'h2b,8'h1a,8'h1b,8'h4,8'h1b,8'h1a,8'h1a,8'h1a,8'h3,8'h21,8'h2b,8'h1a,8'h21,8'h21,8'h1a,8'h1a,8'h1a,8'h2b,8'h1a,8'h21,8'h3,8'h1b,8'h1a,8'h2b,8'h1a,8'h2b,8'h1a,8'h21,8'h21,8'h1a,8'h2b,8'h21,8'h3,8'h1b,8'h21,8'h4,8'h16,8'h1a,8'h21,8'h21,8'h1a,8'h1b,8'h3,8'h1b,8'h2b,8'h2b,8'h1a,8'h1b,8'h3,8'h21,8'h1a,8'h21,8'h21,8'h1a,8'h2b,8'h21,8'h21,8'h1a,8'h21,8'h21,8'h1a,8'h1a,8'h21,8'h21,8'h16,8'h3,8'h21,8'h1a,8'h2b,8'h2b,8'h1a,8'h2b,8'h1a,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h1a,8'h1a,8'h2b,8'h2b,8'h2b,8'h1a,8'h1a,8'h2b,8'h2b,8'h2b,8'h1a,8'h1a,8'h2b,8'h2b,8'h2b,8'h1a,8'h1a,8'h1a,8'h2b,8'h2b,8'h2b,8'h1a,8'h1a,8'h2b,8'h2b,8'h2b,8'h1a,8'h1a,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h1a,8'h1a,8'h1a,8'h1a,8'h1a,8'h2b,8'h1a,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h1a,8'h21,8'h4,8'h1b,8'h2b,8'h2b,8'h1a,8'h2b,8'h1a,8'h21,8'h3,8'h1b,8'h2b,8'h2b,8'h21,8'h3,8'h1b,8'h2b,8'h2b,8'h2b,8'h2b,8'h1a,8'h2b,8'h1a,8'h3,8'h21,8'h1a,8'h1a,8'h2b,8'h1a,8'h21,8'h21,8'h1a,8'h2b,8'h1a,8'h1a,8'h2b,8'h21,8'h21,8'h1a,8'h2b,8'h1a,8'h1a,8'h2b,8'h21,8'h3,8'h1a,8'h2b,8'h21,8'h21,8'h1a,8'h1b,8'h3,8'h21,8'h2b,8'h2b,8'h1a,8'h21,8'h21,8'h16,8'h2b,8'h1a,8'h2b,8'h1a,8'h21,8'h21,8'h1a,8'h1a,8'h2b,8'h2b,8'h1a,8'h1a,8'h1a,8'h1b,8'h4,8'h21,8'h1a,8'h1a,8'h1a,8'h21,8'h3,8'h16,8'h1a,8'h21,8'h21,8'h1a,8'h1a,8'h1a,8'h2b,8'h1a,8'h1b,8'h21,8'h21,8'h16,8'h2b,8'h2b,8'h1a,8'h1a,8'h21,8'h3,8'h1a,8'h1a,8'h3,8'h21,8'h1a,8'h21,8'h3,8'h16,8'h1a,8'h21,8'h21,8'h1a,8'h1b,8'h3,8'h21,8'h1a,8'h2b,8'h1a,8'h1b,8'h4,8'h21,8'h2b,8'h21,8'h3,8'h1b,8'h1a,8'h21,8'h21,8'h2b,8'h21,8'h21,8'h1b,8'h1b,8'h3,8'h21,8'h1a,8'h21,8'h3,8'h1b,8'h2b,8'h1a,8'h1a,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h1a,8'h1a,8'h2b,8'h2b,8'h2b,8'h1a,8'h1a,8'h2b,8'h2b,8'h2b,8'h1a,8'h1a,8'h2b,8'h2b,8'h2b,8'h1a,8'h1a,8'h1a,8'h2b,8'h2b,8'h2b,8'h1a,8'h1a,8'h2b,8'h1a,8'h2b,8'h1a,8'h1a,8'h2b,8'h1a,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h1a,8'h1a,8'h1a,8'h1a,8'h1a,8'h2b,8'h1a,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h21,8'h3,8'h1b,8'h1a,8'h1a,8'h1a,8'h2b,8'h2b,8'h21,8'h21,8'h1a,8'h1a,8'h1a,8'h1a,8'h21,8'h3,8'h3,8'h21,8'h21,8'h1b,8'h21,8'h3,8'h21,8'h21,8'h21,8'h1b,8'h3,8'h3,8'h21,8'h21,8'h1b,8'h1a,8'h2b,8'h2b,8'h2b,8'h1a,8'h21,8'h3,8'h3,8'h21,8'h3,8'h21,8'h1b,8'h21,8'h21,8'h1b,8'h1a,8'h21,8'h21,8'h2b,8'h2b,8'h21,8'h3,8'h21,8'h3,8'h1b,8'h1a,8'h3,8'h2,8'h21,8'h3,8'h21,8'h2b,8'h21,8'h21,8'h1a,8'h1a,8'h2b,8'h2b,8'h2b,8'h2b,8'h1a,8'h1a,8'h21,8'h21,8'h4,8'h4,8'h1b,8'h1a,8'h21,8'h3,8'h3,8'h21,8'h1b,8'h1a,8'h1a,8'h1a,8'h1a,8'h2b,8'h2b,8'h1b,8'h21,8'h21,8'h3,8'h3,8'h21,8'h1b,8'h1b,8'h21,8'h21,8'h3,8'h21,8'h1a,8'h1a,8'h21,8'h21,8'h1a,8'h1a,8'h21,8'h21,8'h1a,8'h1a,8'h21,8'h21,8'h3,8'h3,8'h1b,8'h1b,8'h4,8'h1b,8'h1a,8'h21,8'h3,8'h1a,8'h1a,8'h21,8'h21,8'h2b,8'h1b,8'h21,8'h3,8'h21,8'h3,8'h21,8'h1a,8'h1a,8'h3,8'h3,8'h21,8'h3,8'h21,8'h1a,8'h1a,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h1a,8'h1a,8'h2b,8'h2b,8'h2b,8'h1a,8'h1a,8'h2b,8'h2b,8'h2b,8'h1a,8'h1a,8'h2b,8'h2b,8'h2b,8'h1a,8'h1a,8'h1a,8'h2b,8'h2b,8'h2b,8'h1a,8'h1a,8'h2b,8'h1a,8'h1a,8'h1a,8'h1a,8'h2b,8'h1a,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h1a,8'h1a,8'h1a,8'h1a,8'h1a,8'h2b,8'h1a,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h1a,8'h1a,8'h2b,8'h1a,8'h2b,8'h2b,8'h1a,8'h1a,8'h2b,8'h1a,8'h1a,8'h2b,8'h1a,8'h2b,8'h2b,8'h2b,8'h1a,8'h2b,8'h2b,8'h2b,8'h1a,8'h2b,8'h1a,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h1a,8'h1a,8'h2b,8'h1a,8'h2b,8'h2b,8'h2b,8'h1a,8'h2b,8'h1a,8'h2b,8'h2b,8'h1a,8'h2b,8'h2b,8'h2b,8'h1a,8'h2b,8'h2b,8'h2b,8'h1a,8'h2b,8'h2b,8'h1a,8'h2b,8'h2b,8'h2b,8'h1a,8'h2b,8'h2b,8'h1a,8'h1a,8'h2b,8'h1a,8'h2b,8'h1a,8'h2b,8'h1a,8'h2b,8'h1a,8'h2b,8'h1a,8'h1a,8'h1a,8'h1a,8'h1a,8'h1a,8'h1a,8'h2b,8'h2b,8'h2b,8'h1a,8'h2b,8'h1a,8'h1a,8'h1a,8'h1a,8'h1a,8'h2b,8'h2b,8'h2b,8'h1a,8'h1a,8'h2b,8'h2b,8'h2b,8'h1a,8'h1a,8'h2b,8'h1a,8'h1a,8'h2b,8'h2b,8'h2b,8'h1a,8'h1a,8'h1a,8'h2b,8'h2b,8'h1a,8'h2b,8'h2b,8'h2b,8'h1a,8'h2b,8'h2b,8'h1a,8'h2b,8'h1a,8'h1a,8'h1a,8'h2b,8'h2b,8'h2b,8'h2b,8'h1a,8'h2b,8'h2b,8'h1a,8'h2b,8'h1a,8'h1a,8'h2b,8'h1a,8'h1a,8'h2b,8'h2b,8'h1a,8'h2b,8'h1a,8'h2b,8'h1a,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b};
assign data = screen[addr];

endmodule
