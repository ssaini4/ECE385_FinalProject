module font_pokemon ( input [9:0] addr, output [7:0] data);
					 
parameter ADDR_WIDTH = 10;
parameter DATA_WIDTH = 24;

logic [899:0] addr_reg;

parameter [0:899][DATA_WIDTH-1:0] pokemon_one = {
24'hffffff, 24'hffffff, 24'hffffff, 24'hffffff, 24'hffffff, 24'hffffff, 24'hffffff, 24'hfffcfd, 24'heaffff, 24'hfffbff, 24'hfffbff, 24'hfcffff, 24'hf5fffd, 24'hfff7ff, 24'hf7fffd, 24'hfffdff, 24'hffffff, 24'hffffff, 24'hffffff, 24'hffffff, 24'hffffff, 24'hffffff, 24'hffffff, 24'hffffff, 24'hffffff, 24'hffffff, 24'hffffff, 24'hffffff, 24'hffffff, 24'hffffff, 24'hffffff, 24'hffffff, 24'hffffff, 24'hffffff, 24'hffffff, 24'hffffff, 24'hffffff, 24'hf4ffff, 24'h30aa9f, 24'h5cded2, 24'h78e1e5, 24'h7ae0e2, 24'h2fc1b7, 24'h259191, 24'h357a77, 24'hfffcfa, 24'hffffff, 24'hffffff, 24'hffffff, 24'hffffff, 24'hffffff, 24'hffffff, 24'hffffff, 24'hffffff, 24'hffffff, 24'hffffff, 24'hffffff, 24'hffffff, 24'hffffff, 24'hffffff, 24'hffffff, 24'hffffff, 24'hffffff, 24'hffffff, 24'hffffff, 24'hffffff, 24'hfeffff, 24'h09c8f, 24'h87e7dc, 24'h8de3e4, 24'h8aeeee, 24'h35cad0, 24'h2fceca, 24'h33ccca, 24'h2ccfcc, 24'h16662, 24'hfff9fb, 24'hffffff, 24'hffffff, 24'hffffff, 24'hffffff, 24'hffffff, 24'hffffff, 24'hffffff, 24'hffffff, 24'hffffff, 24'hffffff, 24'hffffff, 24'hffffff, 24'hffffff, 24'hffffff, 24'hffffff, 24'hffffff, 24'hffffff, 24'hffffff, 24'hffffff, 24'h196b67, 24'h83e3df, 24'h7aede0, 24'h87eff0, 24'h30c8c9, 24'h32cccc, 24'h32cccc, 24'h32cccc, 24'h32cccc, 24'h32cccc, 24'hebffff, 24'hfff9f3, 24'hffffff, 24'hffffff, 24'hffffff, 24'hffffff, 24'hffffff, 24'hffffff, 24'hffffff, 24'hffffff, 24'hffffff, 24'hffffff, 24'hffffff, 24'hffffff, 24'hffffff, 24'hffffff, 24'hffffff, 24'hffffff, 24'hffffff, 24'hffffff, 24'h40cacd, 24'h3bc3c3, 24'h2ad0c4, 24'h34cece, 24'h33cbcc, 24'h09696, 24'h32cccc, 24'h32cccc, 24'h32cccc, 24'h32cccc, 24'h8666e, 24'hfdfdfb, 24'hffffff, 24'hffffff, 24'hffffff, 24'hffffff, 24'hffffff, 24'hffffff, 24'hffffff, 24'hffffff, 24'hffffff, 24'hffffff, 24'hffffff, 24'hffffff, 24'hffffff, 24'hffffff, 24'hffffff, 24'hffffff, 24'hfffffa, 24'h26159, 24'h44c6d3, 24'h32cccc, 24'h32cccc, 24'h32cccc, 24'h32cccc, 24'h3bd0d4, 24'h09996, 24'h9929c, 24'h2cd2d0, 24'h2fcec9, 24'h29396, 24'h06a60, 24'hffffff, 24'hffffff, 24'hffffff, 24'hffffff, 24'hffffff, 24'hffffff, 24'hffffff, 24'hffffff, 24'hffffff, 24'hffffff, 24'hffffff, 24'hffffff, 24'hffffff, 24'hffffff, 24'hffffff, 24'hffffff, 24'hfffffa, 24'h06c6e, 24'h51b8b5, 24'h33cdcd, 24'h32cccc, 24'h32cccc, 24'h32cccc, 24'h6757e, 24'h830, 24'hece2ea, 24'h78786, 24'h2fc9c9, 24'h09a9a, 24'h050, 24'hffffff, 24'hffffff, 24'hffffff, 24'hffffff, 24'hffffff, 24'hffffff, 24'hffffff, 24'hffffff, 24'hffffff, 24'hffffff, 24'hffffff, 24'hffffff, 24'hffffff, 24'hffffff, 24'hffffff, 24'hffffff, 24'hf8fffa, 24'h46b67, 24'ha9e7e, 24'h38d0d1, 24'h32cccc, 24'h32cccc, 24'h32cccc, 24'h0c10, 24'h701, 24'hf4e3cf, 24'h06c67, 24'ha959c, 24'h09899, 24'h060, 24'hffffff, 24'hffffff, 24'hffffff, 24'hffffff, 24'hffffff, 24'hffffff, 24'hffffff, 24'hffffff, 24'hffffff, 24'hffffff, 24'hffffff, 24'hffffff, 24'hffffff, 24'hffffff, 24'hffffff, 24'hffffff, 24'hfff2f8, 24'h10646f, 24'h9be6e1, 24'h30caca, 24'h32cccc, 24'h32cccc, 24'h32cccc, 24'he3ffff, 24'h560, 24'hfedfcd, 24'h36566, 24'h09c94, 24'h09899, 24'h060, 24'hffffff, 24'hffffff, 24'hffffff, 24'hffffff, 24'hffffff, 24'hffffff, 24'hffffff, 24'hffffff, 24'hffffff, 24'hffffff, 24'hffffff, 24'hffffff, 24'hffffff, 24'hffffff, 24'hffffff, 24'hffffff, 24'h01212, 24'h8be3e4, 24'h249ea1, 24'h30caca, 24'h1cb6b6, 24'h32cccc, 24'h32cccc, 24'h43ae92, 24'h2fa49e, 24'h43a79d, 24'h09693, 24'h09a97, 24'h09899, 24'h060, 24'hffffff, 24'hffffff, 24'hffffff, 24'hffffff, 24'hffffff, 24'hffffff, 24'hffffff, 24'hffffff, 24'hffffff, 24'hffffff, 24'hffffff, 24'hffffff, 24'hffffff, 24'hf9ffff, 24'hfffaff, 24'hfffdfd, 24'hfff8fe, 24'h126, 24'h45cdcd, 24'h34cccd, 24'h34d0cf, 24'h33ccca, 24'h2ccfcc, 24'h2ececc, 24'h09795, 24'h07175, 24'h09b9d, 24'he919b, 24'h00b, 24'hfbfff4, 24'hfff9ff, 24'h1636e, 24'h06862, 24'h1a5857, 24'hfffcff, 24'hffffff, 24'hffffff, 24'hffffff, 24'hffffff, 24'hffffff, 24'hffffff, 24'hffffff, 24'hffffff, 24'hfefff7, 24'h09f9e, 24'hddffff, 24'hf8ffff, 24'hfff9f9, 24'h030, 24'h3bd0cc, 24'h19b8b4, 24'h36566, 24'h5645c, 24'h26562, 24'h56865, 24'h65354, 24'h0a092, 24'h6959b, 24'h9626a, 24'hfffffd, 24'h5939f, 24'h87e2db, 24'h09da1, 24'h1e8a94, 24'hfffeff, 24'hffffff, 24'hffffff, 24'hffffff, 24'hffffff, 24'hffffff, 24'hffffff, 24'hffffff, 24'hffffff, 24'h1a8b8f, 24'h89e7e7, 24'h87e5e5, 24'h84e6e5, 24'h159191, 24'h01115, 24'h3968c, 24'h685a3f, 24'h60360, 24'h67320, 24'h7f280, 24'hb9ba3, 24'h49898, 24'h0655d, 24'h9a0, 24'h7fe6e3, 24'h91e1e0, 24'h8ee3de, 24'h46665, 24'h2a09f, 24'h000, 24'hffffff, 24'hffffff, 24'hffffff, 24'hffffff, 24'hffffff, 24'hffffff, 24'hffffff, 24'hffffff, 24'hffffff, 24'h26668, 24'h87ebe1, 24'h8ae6e3, 24'h8ae4e5, 24'h8ae4e5, 24'h8ae4e5, 24'h700, 24'h07c92, 24'h1196a7, 24'h09f93, 24'h09f91, 24'h0a191, 24'h40c, 24'hf0d15c, 24'he6d3c2, 24'h8be8ef, 24'h8ae4e2, 24'h82e1e5, 24'h29899, 24'h0d0, 24'hffffff, 24'hffffff, 24'hffffff, 24'hffffff, 24'hffffff, 24'hffffff, 24'hffffff, 24'hffffff, 24'hffffff, 24'hffffff, 24'hfffafb, 24'ha6158, 24'hc8c8d, 24'h78e5e8, 24'h78e5e8, 24'h78e5e8, 24'h0a2a1, 24'h2d6c61, 24'ha102, 24'h1790, 24'h10d0, 24'h1340, 24'hf6c356, 24'hbdcd74, 24'h27067, 24'h8be4e2, 24'h7be7ea, 24'h0989d, 24'h11867e, 24'h0a0, 24'hffffff, 24'hffffff, 24'hffffff, 24'hffffff, 24'hffffff, 24'hffffff, 24'hffffff, 24'hffffff, 24'hffffff, 24'hffffff, 24'hffffff, 24'hffffff, 24'hdfffff, 24'h06669, 24'h0999f, 24'h5969b, 24'hb27d9, 24'he9ad31, 24'hfac751, 24'hb9830, 24'hfccc3c, 24'hffe099, 24'hf4d266, 24'h06c71, 24'h0a185, 24'h29491, 24'h09f9b, 24'h168e8c, 24'h6432d, 24'hfbffff, 24'hfeffff, 24'hfeffff, 24'hfaf9fe, 24'h26668, 24'h06b68, 24'h06b6d, 24'hfffeff, 24'hffffff, 24'hffffff, 24'hffffff, 24'hffffff, 24'hffffff, 24'hfeffff, 24'hfffeff, 24'h700, 24'h050, 24'ha4810, 24'hfbebaf, 24'hb67ce, 24'hecc858, 24'hf7eec3, 24'hf9db93, 24'hf4e195, 24'ha57d4, 24'h06f78, 24'h09b9b, 24'h09d9b, 24'h1340, 24'hb2764, 24'h79390, 24'hf5ffff, 24'h67167, 24'h36564, 24'h8be6e9, 24'h8ad8e2, 24'h29c9c, 24'h176663, 24'hffffff, 24'hffffff, 24'hffffff, 24'hffffff, 24'hffffff, 24'hffffff, 24'hffffff, 24'hffffff, 24'haa81b, 24'hffefc4, 24'hffe9b2, 24'hfac855, 24'hfaebc4, 24'hffecc1, 24'hffecbd, 24'hf2cf73, 24'hf2b443, 24'hfec552, 24'h4b296, 24'hadc1c0, 24'hf2f1ec, 24'hb87c0, 24'h662c0, 24'h3c918e, 24'h64d6d6, 24'h8be4e0, 24'h84dedc, 24'h8bdfe1, 24'h8ae4e4, 24'h59cac8, 24'hf0f8fb, 24'hf9f9f9, 24'hffffff, 24'hffffff, 24'hffffff, 24'hffffff, 24'hffffff, 24'hffffff, 24'had7ff, 24'hfee9bc, 24'hffe9c2, 24'hfac754, 24'hffefc5, 24'hfeedc2, 24'hffebc0, 24'hb58521, 24'hf7dd90, 24'hf3ca4c, 24'h64310, 24'hf1eaf2, 24'hf7f1e5, 24'hbe7818, 24'h09d, 24'h09899, 24'h09899, 24'h91e2e3, 24'h80e0dc, 24'h26668, 24'h88e3de, 24'h6fe3e3, 24'h025, 24'hfffeff, 24'hffffff, 24'hffffff, 24'hffffff, 24'hffffff, 24'hffffff, 24'hffffff, 24'had7ff, 24'hb77d11, 24'hffdaae, 24'hc1808, 24'hffeebf, 24'hfff1b1, 24'hfcda83, 24'hfccb6f, 24'hf1df97, 24'hebca63, 24'hb97d3, 24'hfdebdf, 24'hf9eddf, 24'h400, 24'h64350, 24'h09899, 24'h09899, 24'h59794, 24'h0676a, 24'h8de9e4, 24'h56766, 24'h6ee4e6, 24'h025, 24'hfffeff, 24'hffffff, 24'hffffff, 24'hffffff, 24'hffffff, 24'hffffff, 24'hffffff, 24'hb77e0, 24'hffecd1, 24'hffe8af, 24'hbb778, 24'hfff2b8, 24'hfff1bb, 24'hfee088, 24'hbc88e, 24'hf8dd90, 24'hf7dd90, 24'hbf7a5, 24'h63320, 24'heef7f2, 24'hae808, 24'he00, 24'h09899, 24'h09899, 24'h0f5, 24'h29896, 24'h99a93, 24'h3948d, 24'hc8782, 24'hfbffff, 24'hfffdfe, 24'hffffff, 24'hffffff, 24'hffffff, 24'hffffff, 24'hffffff, 24'hffffff, 24'ha1951d, 24'hf7db7a, 24'hffe8bb, 24'hf3bc55, 24'hfff4d3, 24'hfaf0bb, 24'hfbedca, 24'heecc6b, 24'hb4720, 24'hf7c645, 24'h09aa5, 24'h56563, 24'h77074, 24'ha87fd, 24'hc0d, 24'h09899, 24'h09899, 24'h400, 24'h09d99, 24'h09a97, 24'h09a97, 24'ha817f, 24'hfff9fb, 24'hfffeff, 24'hffffff, 24'hffffff, 24'hffffff, 24'hffffff, 24'he7ffff, 24'h1a8b99, 24'h8ae8cd, 24'hc17d0, 24'hffda71, 24'hf9c74a, 24'hfcd97b, 24'hffe9a0, 24'hffe9a0, 24'hface63, 24'h8b8344, 24'h179ca3, 24'h91e1de, 24'h89e5e0, 24'h169989, 24'hdbfffe, 24'h0f12, 24'h09899, 24'h09899, 24'h0a0a0, 24'h02920, 24'h1c8a81, 24'h1a837c, 24'h0d8, 24'hffffff, 24'hffffff, 24'hffffff, 24'hffffff, 24'hffffff, 24'hffffff, 24'h0a098, 24'h91e6e9, 24'h8ae4e2, 24'h92e4de, 24'hb39f26, 24'hf6c455, 24'hfac752, 24'hbb7b0, 24'hba7a0, 24'hb6780, 24'h06976, 24'h86e2ef, 24'h8ae4e2, 24'h89e5e2, 24'h83e5e4, 24'h065, 24'hc8f99, 24'h09697, 24'h09697, 24'h004, 24'h042, 24'hffffff, 24'hfefefe, 24'hffffff, 24'hffffff, 24'hffffff, 24'hffffff, 24'hffffff, 24'hffffff, 24'hffffff, 24'h116862, 24'h92e0ea, 24'h8ae4e2, 24'h84e7e4, 24'h874a2e, 24'hf3c846, 24'hf4c35a, 24'hf8ca50, 24'hf8ca50, 24'hb87a1, 24'h06269, 24'h76e9f0, 24'h8ae4e2, 24'h87e5e5, 24'h7cefec, 24'h06567, 24'h070, 24'h0c0, 24'h0c0, 24'hfeffff, 24'hfffeff, 24'hffffff, 24'hffffff, 24'hffffff, 24'hffffff, 24'hffffff, 24'hffffff, 24'hffffff, 24'hffffff, 24'hffffff, 24'h807272, 24'h02e24, 24'h25a5a4, 24'h24a6a8, 24'h7988b, 24'h3e6e58, 24'h367546, 24'h7d460, 24'h2c200, 24'h3b1c0, 24'h080, 24'h127282, 24'h29a4a2, 24'h29a3a8, 24'h09899, 24'h09899, 24'h130, 24'hffffff, 24'hffffff, 24'hffffff, 24'hffffff, 24'hffffff, 24'hffffff, 24'hffffff, 24'hffffff, 24'hffffff, 24'hffffff, 24'hffffff, 24'hffffff, 24'hffffff, 24'hfffcf6, 24'h07064, 24'h09997, 24'h09996, 24'h099a4, 24'h0a49b, 24'hc012, 24'hfefcff, 24'hfafbff, 24'hfffff7, 24'hf7fffa, 24'h1d07, 24'he909d, 24'h29897, 24'h09899, 24'h09899, 24'h130, 24'hffffff, 24'hffffff, 24'hffffff, 24'hffffff, 24'hffffff, 24'hffffff, 24'hffffff, 24'hffffff, 24'hffffff, 24'hffffff, 24'hffffff, 24'hffffff, 24'hffffff, 24'h8736d, 24'h80dbd2, 24'h0615d, 24'h85d7d3, 24'h2e5248, 24'h020, 24'hfffeff, 24'hffffff, 24'hffffff, 24'hffffff, 24'hffffff, 24'hffffff, 24'ha9286, 24'h1969a, 24'ha918d, 24'h0a29d, 24'h14959b, 24'h555, 24'hffffff, 24'hffffff, 24'hffffff, 24'hffffff, 24'hffffff, 24'hffffff, 24'hffffff, 24'hffffff, 24'hffffff, 24'hffffff, 24'hffffff, 24'hffffff, 24'hffffff, 24'hffffff, 24'hffffff, 24'hffffff, 24'heeeeee, 24'hffffff, 24'hffffff, 24'hffffff, 24'hffffff, 24'hffffff, 24'hffffff, 24'hffffff, 24'h064, 24'h0e9, 24'hf9ffff, 24'h010d, 24'hfffeff, 24'hffffff, 24'hffffff, 24'hffffff, 24'hffffff, 24'hffffff, 24'hffffff, 24'hffffff, 24'hffffff, 24'hffffff, 24'hffffff, 24'hffffff, 24'hffffff, 24'hffffff, 24'hffffff, 24'hffffff, 24'hffffff, 24'hffffff, 24'hffffff, 24'hffffff, 24'hffffff, 24'hffffff, 24'hffffff, 24'hffffff, 24'hffffff, 24'hffffff, 24'hfffffd, 24'hfffaff, 24'hf8faf9, 24'hfcffff, 24'hfeffff, 24'hffffff, 24'hffffff, 24'hffffff, 24'hffffff, 24'hffffff, 24'hffffff, 24'hffffff, 24'hffffff, 24'hffffff
};
assign data = pokemon_one[addr];

endmodule
