module font_grass ( input [8:0] addr,
					 output [7:0] data
					 );
					 
parameter ADDR_WIDTH = 9;
parameter DATA_WIDTH = 8;

logic [ADDR_WIDTH - 1:0] addr_reg;

parameter [0:400-1][DATA_WIDTH-1:0] grass = {
8'h2,8'h4,8'h4,8'h4,8'h1,8'h4,8'h4,8'h4,8'h4,8'h4,8'h1,8'h4,8'h4,8'h4,8'h2,8'h4,8'h1,8'h4,8'h4,8'h4,8'h4,8'h4,8'h4,8'h1,8'h1,8'h4,8'h1,8'h1,8'h4,8'h1,8'h1,8'h4,8'h4,8'h4,8'h4,8'h1,8'h4,8'h4,8'h1,8'h4,8'h1,8'h1,8'h4,8'h1,8'h4,8'h1,8'h4,8'h2,8'h1,8'h4,8'h4,8'h1,8'h1,8'h4,8'h1,8'h4,8'h4,8'h1,8'h2,8'h4,8'h2,8'h4,8'h4,8'h4,8'h4,8'h1,8'h4,8'h4,8'h4,8'h1,8'h4,8'h2,8'h3,8'h4,8'h4,8'h4,8'h1,8'h4,8'h4,8'h4,8'h4,8'h1,8'h1,8'h4,8'h1,8'h4,8'h4,8'h4,8'h4,8'h4,8'h4,8'h4,8'h1,8'h1,8'h4,8'h4,8'h1,8'h4,8'h4,8'h4,8'h4,8'h4,8'h1,8'h4,8'h4,8'h1,8'h4,8'h1,8'h1,8'h4,8'h4,8'h4,8'h4,8'h1,8'h4,8'h4,8'h1,8'h4,8'h4,8'h1,8'h1,8'h4,8'h3,8'h4,8'h3,8'h1,8'h4,8'h1,8'h4,8'h4,8'h4,8'h1,8'h4,8'h2,8'h4,8'h4,8'h4,8'h1,8'h4,8'h1,8'h1,8'h1,8'h4,8'h4,8'h4,8'h4,8'h4,8'h1,8'h1,8'h1,8'h4,8'h4,8'h1,8'h1,8'h4,8'h4,8'h4,8'h4,8'h4,8'h1,8'h1,8'h0,8'h1,8'h4,8'h4,8'h1,8'h4,8'h1,8'h4,8'h1,8'h1,8'h4,8'h1,8'h0,8'h4,8'h4,8'h4,8'h1,8'h1,8'h1,8'h0,8'h1,8'h1,8'h4,8'h4,8'h4,8'h1,8'h1,8'h1,8'h1,8'h1,8'h0,8'h0,8'h1,8'h4,8'h4,8'h4,8'h1,8'h1,8'h1,8'h0,8'h1,8'h1,8'h4,8'h1,8'h4,8'h4,8'h1,8'h1,8'h1,8'h4,8'h1,8'h0,8'h1,8'h4,8'h1,8'h4,8'h4,8'h1,8'h1,8'h1,8'h3,8'h1,8'h4,8'h3,8'h4,8'h1,8'h1,8'h4,8'h4,8'h1,8'h0,8'h3,8'h1,8'h4,8'h2,8'h4,8'h1,8'h1,8'h4,8'h1,8'h1,8'h1,8'h4,8'h4,8'h1,8'h1,8'h4,8'h4,8'h4,8'h2,8'h1,8'h1,8'h1,8'h4,8'h4,8'h4,8'h1,8'h4,8'h4,8'h4,8'h1,8'h4,8'h2,8'h1,8'h4,8'h4,8'h4,8'h4,8'h4,8'h4,8'h4,8'h1,8'h4,8'h2,8'h4,8'h1,8'h4,8'h3,8'h1,8'h3,8'h4,8'h4,8'h1,8'h1,8'h4,8'h1,8'h1,8'h4,8'h1,8'h1,8'h4,8'h4,8'h4,8'h4,8'h1,8'h4,8'h4,8'h1,8'h4,8'h1,8'h1,8'h4,8'h1,8'h4,8'h4,8'h4,8'h4,8'h1,8'h4,8'h4,8'h1,8'h1,8'h4,8'h4,8'h1,8'h4,8'h1,8'h4,8'h4,8'h3,8'h4,8'h4,8'h1,8'h4,8'h1,8'h4,8'h4,8'h4,8'h1,8'h4,8'h4,8'h4,8'h4,8'h1,8'h4,8'h1,8'h1,8'h4,8'h4,8'h4,8'h4,8'h4,8'h4,8'h1,8'h4,8'h4,8'h4,8'h4,8'h1,8'h4,8'h2,8'h4,8'h1,8'h4,8'h4,8'h1,8'h4,8'h1,8'h2,8'h4,8'h1,8'h1,8'h4,8'h4,8'h1,8'h4,8'h1,8'h1,8'h4,8'h1,8'h4,8'h4,8'h1,8'h4,8'h4,8'h1,8'h4,8'h4,8'h1,8'h4,8'h4,8'h4,8'h4,8'h4,8'h1,8'h4,8'h1,8'h1,8'h4,8'h4,8'h1,8'h4,8'h2,8'h4,8'h4,8'h1,8'h1,8'h4,8'h1};
assign data = grass[addr];

endmodule
