module font_boulder ( input [8:0] addr, input[7:0] keycode,
					 output [7:0] data
					 );
					 
parameter ADDR_WIDTH = 9;
parameter DATA_WIDTH = 8;

parameter [0:400-1][DATA_WIDTH-1:0] boulder = {8'h6,8'h13,8'he,8'h13,8'h10,8'he,8'hc,8'ha,8'ha,8'ha,8'ha,8'hb,8'h13,8'h10,8'h10,8'he,8'he,8'he,8'he,8'h6,8'ha,8'h7,8'h8,8'h12,8'h12,8'h12,8'h12,8'h12,8'h12,8'ha,8'ha,8'hb,8'h10,8'hf,8'h10,8'h10,8'hf,8'h6,8'h6,8'ha,8'h12,8'ha,8'h6,8'h8,8'h7,8'h8,8'h8,8'h7,8'h8,8'h7,8'h7,8'h7,8'h7,8'h7,8'h8,8'h7,8'h8,8'h9,8'h9,8'ha,8'h12,8'h12,8'h7,8'he,8'he,8'h8,8'h11,8'h8,8'h11,8'he,8'h9,8'h8,8'hb,8'h11,8'h8,8'h13,8'ha,8'ha,8'ha,8'ha,8'h12,8'h12,8'h6,8'ha,8'h9,8'ha,8'h8,8'h8,8'h14,8'h9,8'h8,8'h8,8'hb,8'h8,8'hc,8'ha,8'hb,8'ha,8'ha,8'h12,8'h12,8'h12,8'h7,8'h7,8'h12,8'he,8'h11,8'h7,8'h14,8'h8,8'h8,8'h10,8'h7,8'he,8'hb,8'hc,8'h7,8'ha,8'ha,8'h12,8'h12,8'ha,8'h7,8'h10,8'h6,8'hd,8'h13,8'he,8'hf,8'h8,8'h8,8'h8,8'hc,8'hd,8'he,8'h8,8'h8,8'ha,8'ha,8'h12,8'hb,8'ha,8'h7,8'h10,8'h10,8'h6,8'h13,8'hb,8'hd,8'h7,8'h7,8'ha,8'ha,8'h10,8'h6,8'h11,8'h8,8'ha,8'ha,8'ha,8'h12,8'ha,8'h7,8'hf,8'h10,8'h14,8'h8,8'ha,8'ha,8'ha,8'he,8'ha,8'hb,8'h7,8'h10,8'he,8'h8,8'ha,8'ha,8'h12,8'h12,8'hc,8'h7,8'hf,8'hf,8'h14,8'he,8'h6,8'he,8'h10,8'hb,8'ha,8'h7,8'he,8'h10,8'h11,8'h10,8'ha,8'h12,8'h12,8'h12,8'hb,8'h7,8'hf,8'hf,8'h11,8'h11,8'h6,8'h11,8'hb,8'h12,8'ha,8'h8,8'he,8'h10,8'he,8'he,8'hb,8'h12,8'h12,8'h12,8'hd,8'h8,8'h10,8'h10,8'h11,8'h8,8'h10,8'h9,8'hc,8'hb,8'hb,8'hb,8'h7,8'he,8'he,8'he,8'hb,8'h12,8'h12,8'ha,8'hd,8'h8,8'h10,8'h11,8'h8,8'hd,8'ha,8'h13,8'h7,8'h7,8'hc,8'ha,8'ha,8'h7,8'he,8'he,8'hb,8'h12,8'h12,8'ha,8'he,8'h7,8'h10,8'h8,8'hd,8'h12,8'h10,8'h8,8'h11,8'h9,8'h6,8'hc,8'hb,8'ha,8'h8,8'h14,8'he,8'h12,8'h12,8'ha,8'he,8'h17,8'h8,8'h10,8'ha,8'hf,8'h6,8'hc,8'h11,8'h8,8'h8,8'h6,8'he,8'h10,8'h10,8'hf,8'he,8'h12,8'ha,8'h12,8'he,8'h7,8'hd,8'ha,8'h10,8'h7,8'hf,8'h14,8'h14,8'h8,8'h8,8'he,8'h6,8'h10,8'hf,8'ha,8'h9,8'h12,8'hb,8'h12,8'he,8'h8,8'ha,8'h10,8'h8,8'he,8'h9,8'h14,8'h11,8'h8,8'hf,8'he,8'h11,8'h8,8'h13,8'he,8'h9,8'ha,8'he,8'h12,8'h6,8'h9,8'ha,8'ha,8'h12,8'ha,8'ha,8'ha,8'ha,8'ha,8'ha,8'ha,8'ha,8'ha,8'hb,8'h9,8'h6,8'h6,8'hd,8'h12,8'h7,8'h9,8'ha,8'ha,8'ha,8'ha,8'ha,8'ha,8'ha,8'ha,8'ha,8'ha,8'ha,8'h12,8'h12,8'ha,8'hf,8'h6,8'hb,8'h7,8'he,8'he,8'h13,8'h13,8'h13,8'hd,8'ha,8'ha,8'ha,8'ha,8'ha,8'h12,8'ha,8'hb,8'hd,8'he,8'he,8'he,8'h6};
assign data = boulder[addr];
endmodule
