module font_pokeB ( input [9:0] addr, output [7:0] data);
					 
parameter DATA_WIDTH = 8;

parameter [0:899][DATA_WIDTH-1:0] poke = {
8'h2b,8'h2b,8'h2b,8'h2b,8'h21,8'h9,8'h1a,8'h2b,8'h1a,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h1a,8'h1a,8'h2b,8'h1a,8'h1a,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h1a,8'h3,8'h22,8'h21,8'h2b,8'h1a,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h1a,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h1b,8'h9,8'h22,8'h9,8'h1a,8'h2b,8'h1a,8'h1a,8'h1a,8'h2b,8'h1a,8'h1a,8'h1a,8'h2b,8'h2b,8'h1a,8'h1a,8'h21,8'h1b,8'h1a,8'h1a,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h21,8'h6,8'h22,8'hb,8'h16,8'h2b,8'h2b,8'h2b,8'h2b,8'h1a,8'h2b,8'h2b,8'h2b,8'h1a,8'h1b,8'h21,8'h3,8'h9,8'h9,8'h3,8'h1b,8'h2b,8'h1a,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h21,8'h9,8'h9,8'hb,8'h21,8'h2b,8'h1a,8'h1a,8'h1a,8'h2b,8'h2b,8'h16,8'h16,8'h21,8'h9,8'h9,8'h9,8'h2,8'h9,8'h2,8'h1b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h1b,8'ha,8'h20,8'h12,8'ha,8'h16,8'h21,8'h20,8'h20,8'h16,8'h16,8'h20,8'h20,8'h3,8'h9,8'h2,8'h9,8'h9,8'h3,8'h1a,8'h2b,8'h1a,8'h16,8'h1a,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h1a,8'h0,8'h20,8'h20,8'h12,8'h20,8'h18,8'h18,8'h20,8'h20,8'h20,8'h20,8'h1,8'h3,8'h4,8'h9,8'h9,8'h3,8'h1b,8'h2b,8'h2b,8'h16,8'h20,8'h20,8'h1a,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h16,8'h12,8'h20,8'h18,8'h18,8'h18,8'h18,8'h20,8'h20,8'h20,8'h20,8'h20,8'ha,8'h1,8'h21,8'h1b,8'h2b,8'h2b,8'h2b,8'h16,8'h20,8'h20,8'h20,8'h21,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h1b,8'ha,8'h20,8'h20,8'h20,8'h20,8'h20,8'h3,8'h9,8'h0,8'h20,8'ha,8'h21,8'h1a,8'h2b,8'h2b,8'h2b,8'h1a,8'h16,8'h20,8'h20,8'h20,8'h20,8'h20,8'h16,8'h2b,8'h2b,8'h2b,8'h2b,8'h1a,8'ha,8'h9,8'h20,8'h20,8'h20,8'h20,8'h20,8'h9,8'h6,8'h0,8'h20,8'ha,8'h1a,8'h2b,8'h1a,8'h2b,8'h1a,8'h20,8'h20,8'h20,8'h20,8'h20,8'h20,8'h20,8'h1b,8'h2b,8'h2b,8'h2b,8'h2b,8'h1a,8'h1,8'h9,8'h20,8'h20,8'h20,8'h20,8'h20,8'h0,8'h0,8'h20,8'h20,8'h20,8'h21,8'h1a,8'h2b,8'h1a,8'h20,8'h20,8'h20,8'h20,8'h20,8'h20,8'h20,8'h20,8'h20,8'h2b,8'h2b,8'h2b,8'h2b,8'h1b,8'h12,8'h20,8'h20,8'h12,8'h12,8'h12,8'h20,8'h20,8'h20,8'h12,8'h12,8'h12,8'h4,8'h2b,8'h1a,8'h20,8'h20,8'h20,8'h20,8'h20,8'h20,8'h20,8'h20,8'h20,8'h12,8'h2b,8'h2b,8'h2b,8'h2b,8'h21,8'h12,8'h20,8'h20,8'h12,8'h11,8'h1d,8'h12,8'h20,8'h20,8'h1d,8'h1d,8'h12,8'h4,8'h2b,8'h16,8'h20,8'h20,8'h20,8'h20,8'h20,8'h20,8'h20,8'h20,8'h0,8'h21,8'h2b,8'h2b,8'h2b,8'h2b,8'h1b,8'ha,8'h20,8'h20,8'h20,8'h12,8'ha,8'h12,8'h20,8'h20,8'h12,8'h12,8'h24,8'h3,8'h16,8'h20,8'h20,8'h20,8'h20,8'h20,8'h20,8'h20,8'h20,8'h0,8'h21,8'h1a,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h1b,8'ha,8'h20,8'h20,8'h24,8'h12,8'h12,8'h20,8'h20,8'h20,8'h20,8'h20,8'h9,8'ha,8'h20,8'h20,8'h20,8'h20,8'h20,8'h20,8'h0,8'h4,8'h21,8'h1a,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h1a,8'hb,8'h20,8'h20,8'h20,8'h20,8'h20,8'h20,8'h20,8'h20,8'h20,8'h20,8'h0,8'h21,8'h20,8'h20,8'h20,8'h20,8'h12,8'ha,8'h21,8'h1a,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h16,8'h4,8'h20,8'h20,8'h20,8'h20,8'h20,8'h20,8'h20,8'h20,8'h20,8'h20,8'h0,8'h1b,8'h1a,8'h20,8'h20,8'h12,8'h21,8'h1a,8'h2b,8'h2b,8'h2b,8'h1a,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h1b,8'hb,8'h20,8'h20,8'h20,8'h20,8'h20,8'h20,8'h20,8'h20,8'h20,8'h20,8'h0,8'h21,8'h2b,8'h21,8'h12,8'h20,8'h1b,8'h2b,8'h2b,8'h1a,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h1a,8'h21,8'h0,8'h20,8'h20,8'h20,8'h20,8'h20,8'h20,8'h20,8'h20,8'h20,8'h20,8'h0,8'h3,8'h21,8'ha,8'h20,8'h20,8'ha,8'h1b,8'h2b,8'h1a,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h1a,8'h3,8'h20,8'h20,8'h20,8'h20,8'h20,8'h20,8'h20,8'h20,8'h20,8'h20,8'h20,8'h20,8'h9,8'ha,8'h24,8'h20,8'ha,8'ha,8'h1b,8'h2b,8'h1a,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h1a,8'h3,8'h20,8'h20,8'h20,8'h20,8'h20,8'h12,8'h20,8'h20,8'h20,8'h24,8'h20,8'h20,8'h9,8'hc,8'h24,8'h20,8'h1b,8'h16,8'h2b,8'h1a,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h3,8'h12,8'h20,8'h20,8'h20,8'h20,8'ha,8'h12,8'h20,8'h20,8'h20,8'h20,8'h20,8'hb,8'h9,8'hb,8'ha,8'h1a,8'h2b,8'h1a,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h21,8'h0,8'h20,8'h20,8'h20,8'h20,8'h20,8'h20,8'h12,8'h12,8'h20,8'h20,8'h20,8'h20,8'h24,8'h9,8'hb,8'h13,8'ha,8'h1a,8'h2b,8'h1a,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h17,8'h20,8'h20,8'h20,8'h20,8'h20,8'h20,8'h20,8'h20,8'h20,8'h20,8'h20,8'h20,8'h20,8'h20,8'h9,8'h9,8'h9,8'h21,8'h1a,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h23,8'h20,8'h20,8'h20,8'h20,8'h20,8'h20,8'h20,8'h20,8'h20,8'h20,8'h20,8'h20,8'h20,8'h20,8'h12,8'h3,8'h1b,8'h1a,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'ha,8'h20,8'h20,8'h20,8'h20,8'h20,8'h20,8'h20,8'h20,8'h20,8'h20,8'h20,8'h20,8'h20,8'h20,8'h20,8'h1a,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h16,8'ha,8'h24,8'h20,8'h20,8'h24,8'h12,8'ha,8'h12,8'h20,8'h20,8'h20,8'h20,8'h20,8'h12,8'h21,8'h2b,8'h1a,8'h1a,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h1b,8'hb,8'h12,8'h12,8'h12,8'hb,8'h21,8'h21,8'h21,8'ha,8'hb,8'h12,8'h20,8'h12,8'h3,8'h1a,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h1,8'hb,8'ha,8'ha,8'h3,8'h1b,8'h2b,8'h2b,8'h2b,8'h1b,8'h9,8'h9,8'h20,8'h12,8'ha,8'h1a,8'h2b,8'h1a,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h16,8'h21,8'h21,8'h1a,8'h1a,8'h2b,8'h2b,8'h1a,8'h2b,8'h2b,8'h1a,8'h21,8'h3,8'h9,8'h21,8'h1a,8'h2b,8'h1a,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b
};
assign data = poke[addr];

endmodule
