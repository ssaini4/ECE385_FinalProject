module font_rock ( input [9:0] addr, output [7:0] data);
					 
parameter DATA_WIDTH = 8;

parameter [0:399][DATA_WIDTH-1:0] rock = {8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h8,8'h8,8'hf,8'h11,8'h10,8'h7,8'h2b,8'h2b,8'h2b,8'h1c,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'hf,8'h1d,8'h1d,8'h1d,8'h15,8'h1d,8'h15,8'h1d,8'h10,8'h2b,8'h2b,8'h1c,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h5,8'h2b,8'h2b,8'h11,8'h1d,8'h12,8'h12,8'h12,8'h12,8'h15,8'h15,8'h15,8'h11,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h8,8'h2b,8'h8,8'h8,8'hf,8'h11,8'h12,8'h12,8'h12,8'h20,8'h20,8'h20,8'h20,8'h12,8'hc,8'h2b,8'h2b,8'h2b,8'h2b,8'h7,8'h5,8'h2b,8'h10,8'h11,8'hf,8'h1d,8'h12,8'h12,8'h20,8'h20,8'h12,8'h15,8'h20,8'h20,8'hc,8'h10,8'h10,8'h2b,8'h2b,8'h1c,8'h8,8'h2b,8'h11,8'h10,8'h12,8'h20,8'h20,8'h12,8'h12,8'h15,8'h15,8'h15,8'h12,8'h12,8'h10,8'h11,8'h15,8'h13,8'h2b,8'h2b,8'h2b,8'h8,8'hf,8'h10,8'h12,8'h12,8'h20,8'h20,8'h15,8'h15,8'h15,8'h15,8'h15,8'h15,8'h11,8'h1d,8'h20,8'ha,8'h2b,8'h2b,8'h7,8'h11,8'hf,8'h10,8'h11,8'h1d,8'h1d,8'h12,8'h12,8'h15,8'h20,8'h20,8'h12,8'h15,8'h15,8'h1d,8'h12,8'h1d,8'hf,8'h2b,8'h12,8'h15,8'h11,8'h10,8'h11,8'h11,8'h11,8'h1d,8'h11,8'h12,8'h12,8'h1e,8'h20,8'h12,8'h1d,8'h11,8'h1d,8'h1e,8'h9,8'h2b,8'h12,8'h15,8'h11,8'h8,8'hf,8'h11,8'h10,8'h11,8'h11,8'h1d,8'h12,8'h1d,8'h12,8'h11,8'h10,8'h10,8'h1d,8'h12,8'h9,8'h2b,8'hf,8'h11,8'h11,8'hf,8'hf,8'h10,8'h10,8'h10,8'h11,8'h12,8'h12,8'h12,8'h11,8'h11,8'h8,8'h2b,8'h10,8'hf,8'h7,8'h2b,8'h7,8'h10,8'h10,8'h11,8'h11,8'hf,8'hf,8'h10,8'h11,8'h1d,8'h12,8'h11,8'h11,8'h11,8'h8,8'hf,8'h11,8'hf,8'h2b,8'h2b,8'h2b,8'h2b,8'h8,8'h1d,8'h11,8'h10,8'h10,8'h10,8'h10,8'h11,8'h11,8'h11,8'h11,8'h1d,8'h11,8'hc,8'h12,8'hf,8'h2b,8'h2b,8'h2b,8'h2b,8'hf,8'h10,8'h10,8'h10,8'h10,8'hf,8'h10,8'h11,8'h11,8'ha,8'h1d,8'h20,8'h12,8'h11,8'h12,8'h2b,8'h2b,8'h1c,8'h2b,8'h7,8'h11,8'hf,8'hf,8'h8,8'hf,8'h10,8'h11,8'h1d,8'h1d,8'h15,8'h15,8'h12,8'h11,8'h8,8'h7,8'h2b,8'h23,8'h2b,8'h5,8'h2b,8'hf,8'h11,8'h10,8'h2b,8'h2b,8'h10,8'h11,8'h11,8'h1d,8'h12,8'h12,8'h12,8'h1d,8'hf,8'h2b,8'h2b,8'h2b,8'h2b,8'h5,8'h2b,8'h7,8'h11,8'h11,8'h11,8'hf,8'hf,8'hf,8'hf,8'h11,8'h11,8'h11,8'h11,8'hf,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h8,8'h11,8'h11,8'hf,8'h10,8'hf,8'hf,8'hf,8'h10,8'hf,8'h2b,8'h2b,8'h2b,8'h7,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h8,8'hf,8'h10,8'h11,8'h11,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h2b,8'h8,8'h7,8'h7,8'h7,8'h2b,8'h13,8'h5,8'h2b,8'h2b,8'h2b,8'h2b
};
assign data = rock[addr];

endmodule
