module font_player_image ( input [8:0] addr, input[7:0] keycode,
					 output [23:0] data
					 );
					 
parameter ADDR_WIDTH = 9;
parameter DATA_WIDTH = 24;

logic [ADDR_WIDTH - 1:0] addr_reg;
logic [DATA_WIDTH-1:0] temp;
parameter [0:281-1][DATA_WIDTH-1:0] player_sit = {24'hff260, 24'hff260, 24'hff260, 24'hff260, 24'h882840, 24'h882840, 24'h882840, 24'h882840, 24'h882840, 24'h882840, 24'hff260, 24'hff260, 24'hff260, 24'hff260, 24'hff260, 24'hff260, 24'h000, 24'h882840, 24'hf06848, 24'hf06848, 24'hf06848, 24'hf06848, 24'hf06848, 24'hf06848, 24'h882840, 24'h000, 24'hff260, 24'hff260, 24'hff260, 24'hff260, 24'hc03838, 24'hf06848, 24'hf06848, 24'hf06848, 24'hf06848, 24'hf06848, 24'hf06848, 24'hf06848, 24'hf06848, 24'hc03838, 24'hff260, 24'hff260, 24'hff260, 24'hff260, 24'hf06848, 24'hf06848, 24'hf06848, 24'hf06848, 24'hf06848, 24'hf06848, 24'hf06848, 24'hf06848, 24'hf06848, 24'hf06848, 24'hff260, 24'hff260, 24'hff260, 24'h000, 24'hf06848, 24'hf06848, 24'hf06848, 24'hf06848, 24'hf06848, 24'hf06848, 24'hf06848, 24'hf06848, 24'hf06848, 24'hf06848, 24'h000, 24'hff260, 24'hff260, 24'h000, 24'hf06848, 24'hf06848, 24'hf06848, 24'hf06848, 24'hf06848, 24'hf06848, 24'hf06848, 24'hf06848, 24'hf06848, 24'hf06848, 24'h000, 24'hff260, 24'hff260, 24'h000, 24'hc03838, 24'hf06848, 24'hf06848, 24'hf06848, 24'hf06848, 24'hf06848, 24'hf06848, 24'hf06848, 24'hf06848, 24'hc03838, 24'h000, 24'hff260, 24'hff260, 24'h000, 24'hc03838, 24'hc03838, 24'hc03838, 24'hf06848, 24'hf06848, 24'hf06848, 24'hf06848, 24'hc03838, 24'hc03838, 24'hc03838, 24'h000, 24'hff260, 24'hff260, 24'h882840, 24'hc03838, 24'hc03838, 24'hc03838, 24'hc03838, 24'he8e8f8, 24'he8e8f8, 24'hc03838, 24'hc03838, 24'hc03838, 24'hc03838, 24'h882840, 24'hff260, 24'h503018, 24'h503018, 24'hb8b0d0, 24'hc03838, 24'hc03838, 24'hb8b0d0, 24'hc03838, 24'hc03838, 24'hb8b0d0, 24'hc03838, 24'hc03838, 24'hb8b0d0, 24'h503018, 24'h503018, 24'h784040, 24'hd8a078, 24'h503018, 24'h000, 24'hb8b0d0, 24'hb8b0d0, 24'hb8b0d0, 24'hb8b0d0, 24'hb8b0d0, 24'hb8b0d0, 24'h000, 24'h503018, 24'hd8a078, 24'h784040, 24'hff260, 24'h000, 24'h885028, 24'h503018, 24'h384040, 24'h000, 24'h000, 24'h000, 24'h000, 24'h384040, 24'h503018, 24'h885028, 24'h000, 24'hff260, 24'hff260, 24'hff260, 24'hd8a078, 24'hd8a078, 24'hb8b0d0, 24'h000, 24'h784040, 24'h784040, 24'h000, 24'hb8b0d0, 24'hd8a078, 24'hd8a078, 24'hff260, 24'hff260, 24'hff260, 24'hff260, 24'h784040, 24'h784040, 24'hf8d0b8, 24'hf8d0b8, 24'hf8d0b8, 24'hf8d0b8, 24'hf8d0b8, 24'hf8d0b8, 24'h784040, 24'h784040, 24'hff260, 24'hff260, 24'hff260, 24'h000, 24'hf8d0b8, 24'h885028, 24'h000, 24'h784040, 24'hd8a078, 24'hd8a078, 24'h784040, 24'h000, 24'h885028, 24'hf8d0b8, 24'h000, 24'hff260, 24'hff260, 24'h000, 24'hd8a078, 24'h885028, 24'hc03838, 24'hb8b0d0, 24'h784040, 24'h784040, 24'hb8b0d0, 24'hc03838, 24'h885028, 24'hd8a078, 24'h000, 24'hff260, 24'hff260, 24'hff260, 24'h000, 24'h000, 24'hc03838, 24'hc03838, 24'hb8b0d0, 24'hb8b0d0, 24'hc03838, 24'hc03838, 24'h000, 24'h000, 24'hff260, 24'hff260, 24'hff260, 24'hff260, 24'h000, 24'h406888, 24'h384040, 24'hc03838, 24'hb8b0d0, 24'hb8b0d0, 24'hc03838, 24'h384040, 24'h406888, 24'h000, 24'hff260, 24'hff260, 24'hff260, 24'hff260, 24'h000, 24'hc03838, 24'hc03838, 24'h000, 24'h384040, 24'h384040, 24'h000, 24'hc03838, 24'hc03838, 24'h000, 24'hff260, 24'hff260, 24'hff260, 24'hff260, 24'hff260, 24'h000, 24'h000, 24'hff260, 24'hff260, 24'hff260, 24'hff260, 24'h000, 24'h000, 24'hff260, 24'hff260, 24'hff260};
parameter [0:281-1][DATA_WIDTH-1:0] player_walkup = {24'hff9191, 24'hff2626, 24'hff00, 24'hff00, 24'h882840, 24'h882840, 24'h882840, 24'h882840, 24'h882840, 24'h882840, 24'hff00, 24'hff00, 24'hff2626, 24'hff9191, 24'hff2626, 24'hff00, 24'h000, 24'h882840, 24'hf06848, 24'hf06848, 24'hf06848, 24'hf06848, 24'hf06848, 24'hf06848, 24'h882840, 24'h000, 24'hff00, 24'hff2626, 24'hff00, 24'hff00, 24'hf06848, 24'hf06848, 24'hf06848, 24'hf06848, 24'hf06848, 24'hf06848, 24'hf06848, 24'hf06848, 24'hf06848, 24'hf06848, 24'hff00, 24'hff00, 24'hff00, 24'h000, 24'hf06848, 24'hf06848, 24'hf06848, 24'hf06848, 24'hf06848, 24'hf06848, 24'hf06848, 24'hf06848, 24'hf06848, 24'hf06848, 24'h000, 24'hff00, 24'hff00, 24'h000, 24'hf06848, 24'hf06848, 24'hf06848, 24'hf06848, 24'hf06848, 24'hf06848, 24'hf06848, 24'hf06848, 24'hf06848, 24'hf06848, 24'h000, 24'hff00, 24'hff00, 24'h000, 24'hc03838, 24'hf06848, 24'hf06848, 24'hf06848, 24'hf06848, 24'hf06848, 24'hf06848, 24'hf06848, 24'hf06848, 24'hc03838, 24'h000, 24'hff00, 24'h503018, 24'h882840, 24'hc03838, 24'hc03838, 24'hc03838, 24'hc03838, 24'h384040, 24'h384040, 24'hc03838, 24'hc03838, 24'hc03838, 24'hc03838, 24'h882840, 24'hff00, 24'h000, 24'hd8a078, 24'hc03838, 24'hc03838, 24'hc03838, 24'h384040, 24'h384040, 24'h384040, 24'h384040, 24'hc03838, 24'hc03838, 24'hc03838, 24'hd8a078, 24'h000, 24'h000, 24'hd8a078, 24'h000, 24'h000, 24'hc03838, 24'hc03838, 24'hc03838, 24'hc03838, 24'hc03838, 24'hc03838, 24'h000, 24'h000, 24'hd8a078, 24'h000, 24'hff00, 24'h000, 24'h885028, 24'h503018, 24'h000, 24'h000, 24'h000, 24'h000, 24'h000, 24'h000, 24'h503018, 24'h885028, 24'h000, 24'hff00, 24'h000, 24'hd8a078, 24'h000, 24'h503018, 24'h885028, 24'h885028, 24'h885028, 24'h885028, 24'h885028, 24'h885028, 24'h503018, 24'h000, 24'hff00, 24'hff00, 24'hff00, 24'h000, 24'h384040, 24'h000, 24'h000, 24'h503018, 24'h885028, 24'h885028, 24'h503018, 24'h000, 24'h000, 24'hff00, 24'hff00, 24'hff00, 24'hff00, 24'hff00, 24'h384040, 24'h882840, 24'hc8980, 24'h503018, 24'h503018, 24'h503018, 24'h503018, 24'hc8980, 24'h384040, 24'h000, 24'hff00, 24'hff00, 24'hff00, 24'hff00, 24'h000, 24'hc03838, 24'h000, 24'h885028, 24'hc8980, 24'hc8980, 24'h885028, 24'h000, 24'h384040, 24'h000, 24'hff00, 24'hff00, 24'hff00, 24'hff00, 24'h406888, 24'h000, 24'h503018, 24'hc8980, 24'hc8980, 24'hc8980, 24'hc8980, 24'h503018, 24'h000, 24'h000, 24'hff00, 24'hff00, 24'hff00, 24'hff00, 24'h000, 24'h406888, 24'h406888, 24'h000, 24'hc8980, 24'hc8980, 24'h000, 24'h384040, 24'h384040, 24'hf8d0b8, 24'h000, 24'hff00, 24'hff00, 24'hff00, 24'h000, 24'h406888, 24'h406888, 24'h000, 24'h000, 24'h406888, 24'h384040, 24'h000, 24'h406888, 24'hd8a078, 24'h000, 24'hff00, 24'hff00, 24'hff00, 24'h000, 24'h406888, 24'h406888, 24'h384040, 24'h000, 24'h000, 24'hff00, 24'hff00, 24'hff00, 24'h000, 24'hff00, 24'hff00, 24'hff2626, 24'hff00, 24'hff00, 24'h000, 24'hf06848, 24'hf06848, 24'h000, 24'hff00, 24'hff00, 24'hff00, 24'hff00, 24'hff00, 24'hff00, 24'hff2626, 24'hff9191, 24'hff2626, 24'hff00, 24'hff00, 24'h000, 24'h000, 24'hff00, 24'hff00, 24'hff00, 24'hff00, 24'hff00, 24'hff00, 24'hff2626, 24'hff9191};
parameter [0:281-1][DATA_WIDTH-1:0] player_walkright = {24'hff9191, 24'hff2626, 24'hff00, 24'hff00, 24'h882840, 24'h882840, 24'h882840, 24'h882840, 24'h882840, 24'h882840, 24'hff00, 24'hff00, 24'hff2626, 24'hff9191, 24'hff2626, 24'hff00, 24'h000, 24'h882840, 24'hf06848, 24'hf06848, 24'hf06848, 24'hf06848, 24'hf06848, 24'hc03838, 24'h882840, 24'hff00, 24'hff00, 24'hff2626, 24'hff00, 24'hff00, 24'hc03838, 24'hf06848, 24'hf06848, 24'hf06848, 24'hf06848, 24'hf06848, 24'hf06848, 24'hf06848, 24'hc03838, 24'h882840, 24'hff00, 24'hff00, 24'hff00, 24'h882840, 24'hf06848, 24'hf06848, 24'hf06848, 24'hf06848, 24'hf06848, 24'hf06848, 24'hf06848, 24'hf06848, 24'hf06848, 24'hb8b0d0, 24'hff00, 24'hff00, 24'hff00, 24'h000, 24'hf06848, 24'hf06848, 24'hf06848, 24'hf06848, 24'hf06848, 24'hf06848, 24'hf06848, 24'hf06848, 24'he8e8f8, 24'hc03838, 24'h384040, 24'hff00, 24'hff00, 24'h000, 24'hc03838, 24'hf06848, 24'hf06848, 24'hf06848, 24'hf06848, 24'hf06848, 24'hf06848, 24'hc03838, 24'he8e8f8, 24'hc03838, 24'he8e8f8, 24'h000, 24'hff00, 24'h000, 24'hc03838, 24'hc03838, 24'hc03838, 24'hc03838, 24'hc03838, 24'hc03838, 24'hc03838, 24'hc03838, 24'hc03838, 24'hb8b0d0, 24'he8e8f8, 24'h000, 24'hff00, 24'h000, 24'hc03838, 24'hc03838, 24'hc03838, 24'hc03838, 24'hc03838, 24'hc03838, 24'hc03838, 24'hc03838, 24'hc03838, 24'h882840, 24'hb8b0d0, 24'h000, 24'hff00, 24'h503018, 24'hc03838, 24'hc03838, 24'hc03838, 24'hc03838, 24'hc03838, 24'hc03838, 24'hc03838, 24'hc03838, 24'h882840, 24'hb8b0d0, 24'h000, 24'hff00, 24'hff00, 24'h503018, 24'h000, 24'h000, 24'h000, 24'h000, 24'h000, 24'h000, 24'h000, 24'h000, 24'h384040, 24'h000, 24'hff00, 24'hff00, 24'hff00, 24'hff00, 24'h503018, 24'h885028, 24'h885028, 24'h503018, 24'hd8a078, 24'h503018, 24'hd8a078, 24'he8e8f8, 24'h000, 24'hd8a078, 24'hff00, 24'hff00, 24'hff00, 24'hff00, 24'h000, 24'h885028, 24'h885028, 24'h503018, 24'hd8a078, 24'hd8a078, 24'hf8d0b8, 24'hf8d0b8, 24'hf8d0b8, 24'hf8d0b8, 24'hff00, 24'hff00, 24'hff00, 24'h503018, 24'h503018, 24'h503018, 24'h000, 24'h503018, 24'h503018, 24'hd8a078, 24'hd8a078, 24'hf8d0b8, 24'hf8d0b8, 24'h784040, 24'hff00, 24'hff00, 24'h503018, 24'hc8980, 24'hc8980, 24'h885028, 24'h885028, 24'hc8980, 24'h885028, 24'h000, 24'h784040, 24'h784040, 24'h784040, 24'hff00, 24'hff00, 24'hff00, 24'h000, 24'h885028, 24'hc8980, 24'h000, 24'hc03838, 24'hc03838, 24'h882840, 24'h384040, 24'h000, 24'h000, 24'hff00, 24'hff00, 24'hff00, 24'hff00, 24'h000, 24'hc8980, 24'h000, 24'hc03838, 24'hc03838, 24'hc03838, 24'h000, 24'h000, 24'hf8d0b8, 24'hf8d0b8, 24'h784040, 24'hff00, 24'hff00, 24'hff00, 24'h000, 24'h885028, 24'h000, 24'h784040, 24'hc03838, 24'hc03838, 24'hc03838, 24'h000, 24'hd8a078, 24'hd8a078, 24'h784040, 24'hff00, 24'hff00, 24'hff00, 24'h000, 24'hc03838, 24'h406888, 24'h406888, 24'h406888, 24'h406888, 24'h000, 24'h384040, 24'h384040, 24'hc03838, 24'h000, 24'hff00, 24'hff00, 24'hff00, 24'h000, 24'hc03838, 24'h000, 24'h000, 24'h000, 24'h000, 24'hff00, 24'hff00, 24'h000, 24'h000, 24'hff00, 24'hff00, 24'hff00, 24'hff2626, 24'hff9191, 24'h000, 24'hff00, 24'hff00, 24'hff00, 24'hff00, 24'hff00, 24'hff00, 24'hff00, 24'hff00, 24'hff00, 24'hff00, 24'hff2626, 24'hff9191};
parameter [0:281-1][DATA_WIDTH-1:0] player_walkleft = {24'hff9191, 24'hff2626, 24'hff00, 24'hff00, 24'h882840, 24'h882840, 24'h882840, 24'h882840, 24'h882840, 24'h882840, 24'hff00, 24'hff00, 24'hff2525, 24'hff9191, 24'hff2626, 24'hff00, 24'hff00, 24'h882840, 24'hc03838, 24'hf06848, 24'hf06848, 24'hf06848, 24'hf06848, 24'hf06848, 24'h882840, 24'h400, 24'hff00, 24'hff2121, 24'hff00, 24'hff00, 24'h882840, 24'hc03838, 24'hf06848, 24'hf06848, 24'hf06848, 24'hf06848, 24'hf06848, 24'hf06848, 24'hf06848, 24'hc03838, 24'hff00, 24'hff00, 24'hff00, 24'hff00, 24'hb8b0d0, 24'hf06848, 24'hf06848, 24'hf06848, 24'hf06848, 24'hf06848, 24'hf06848, 24'hf06848, 24'hf06848, 24'hf06848, 24'h8c273e, 24'hff00, 24'hff00, 24'h384040, 24'hc03838, 24'he8e8f8, 24'hf06848, 24'hf06848, 24'hf06848, 24'hf06848, 24'hf06848, 24'hf06848, 24'hf06848, 24'hf06848, 24'h000, 24'hff00, 24'h000, 24'he8e8f8, 24'hc03838, 24'he8e8f8, 24'hc03838, 24'hf06848, 24'hf06848, 24'hf06848, 24'hf06848, 24'hf06848, 24'hf06848, 24'hc03838, 24'h000, 24'hff00, 24'h000, 24'he8e8f8, 24'hb8b0d0, 24'hc03838, 24'hc03838, 24'hc03838, 24'hc03838, 24'hc03838, 24'hc03838, 24'hc03838, 24'hc03838, 24'hc03838, 24'h000, 24'hff00, 24'h000, 24'hb8b0d0, 24'h882840, 24'hc03838, 24'hc03838, 24'hc03838, 24'hc03838, 24'hc03838, 24'hc03838, 24'hc03838, 24'hc03838, 24'hc03838, 24'h000, 24'hff00, 24'hff00, 24'h000, 24'hb8b0d0, 24'h882840, 24'hc03838, 24'hc03838, 24'hc03838, 24'hc03838, 24'hc03838, 24'hc03838, 24'hc03838, 24'hc03838, 24'h503018, 24'hff00, 24'hff00, 24'hff00, 24'h000, 24'h384040, 24'h000, 24'h000, 24'h000, 24'h000, 24'h000, 24'h000, 24'h000, 24'h000, 24'h503018, 24'hff00, 24'hff00, 24'hff00, 24'hd8a078, 24'h000, 24'he8e8f8, 24'hd8a078, 24'h503018, 24'hd8a078, 24'h503018, 24'h885028, 24'h885028, 24'h503018, 24'hff00, 24'hff00, 24'hff00, 24'hff00, 24'hf8d0b8, 24'hf8d0b8, 24'hf8d0b8, 24'hf8d0b8, 24'hd8a078, 24'hd8a078, 24'h503018, 24'h885028, 24'h885028, 24'h000, 24'hff00, 24'hff00, 24'hff00, 24'hff00, 24'h784040, 24'hf8d0b8, 24'hf8d0b8, 24'hd8a078, 24'hd8a078, 24'h503018, 24'h503018, 24'h000, 24'h503018, 24'h503018, 24'h503018, 24'hff00, 24'hff00, 24'hff00, 24'hff00, 24'h784040, 24'h784040, 24'h784040, 24'h000, 24'h885028, 24'hc8980, 24'h885028, 24'h885028, 24'hc8980, 24'hc8980, 24'h503018, 24'hff00, 24'hff00, 24'hff00, 24'hff00, 24'h000, 24'h000, 24'h384040, 24'h882840, 24'hc03838, 24'hc03838, 24'h000, 24'hc8980, 24'h885028, 24'h000, 24'hff00, 24'hff00, 24'hff00, 24'h784040, 24'hf8d0b8, 24'hf8d0b8, 24'h000, 24'h000, 24'hc03838, 24'hc03838, 24'hc03838, 24'h000, 24'hc8980, 24'h000, 24'hff00, 24'hff00, 24'hff00, 24'h784040, 24'hd8a078, 24'hd8a078, 24'h000, 24'hc03838, 24'hc03838, 24'hc03838, 24'h784040, 24'h000, 24'h885028, 24'h000, 24'hff00, 24'hff00, 24'hff00, 24'h000, 24'hc03838, 24'h384040, 24'h384040, 24'h000, 24'h406888, 24'h406888, 24'h406888, 24'h406888, 24'hc03838, 24'h000, 24'hff2626, 24'hff00, 24'hff00, 24'hff00, 24'h000, 24'h000, 24'hff00, 24'hff00, 24'h000, 24'h000, 24'h000, 24'h000, 24'hc03838, 24'h000, 24'hff9191, 24'hff2626, 24'hff00, 24'hff00, 24'hff00, 24'hff00, 24'hff00, 24'hff00, 24'hff00, 24'hff00, 24'hff00, 24'hff00, 24'h000, 24'hff9191};
parameter [0:281-1][DATA_WIDTH-1:0] player_walkdown = {24'hff9191, 24'hff2626, 24'hff00, 24'h882840, 24'h882840, 24'h882840, 24'h882840, 24'h882840, 24'hff00, 24'hff00, 24'hff00, 24'hff00, 24'hff2626, 24'hff9191, 24'hff2626, 24'hff00, 24'h000, 24'hf06848, 24'hf06848, 24'hf06848, 24'hf06848, 24'hf06848, 24'h882840, 24'h000, 24'hff00, 24'hff00, 24'hff00, 24'hff2626, 24'hff00, 24'h000, 24'hc03838, 24'hf06848, 24'hf06848, 24'hf06848, 24'hf06848, 24'hf06848, 24'hf06848, 24'hc03838, 24'hff00, 24'hff00, 24'hff00, 24'hff00, 24'hff00, 24'hc03838, 24'hf06848, 24'hf06848, 24'hf06848, 24'hf06848, 24'hf06848, 24'hf06848, 24'hf06848, 24'hf06848, 24'h000, 24'hff00, 24'hff00, 24'hff00, 24'hff00, 24'hc03838, 24'hf06848, 24'hf06848, 24'hf06848, 24'hf06848, 24'hf06848, 24'hf06848, 24'hf06848, 24'hf06848, 24'h000, 24'hff00, 24'hff00, 24'hff00, 24'hff00, 24'hc03838, 24'hc03838, 24'hf06848, 24'hf06848, 24'hf06848, 24'hf06848, 24'hf06848, 24'hf06848, 24'hc03838, 24'h000, 24'hff00, 24'hff00, 24'hff00, 24'hff00, 24'hc03838, 24'hc03838, 24'hc03838, 24'hf06848, 24'hf06848, 24'hf06848, 24'hf06848, 24'hc03838, 24'hc03838, 24'h000, 24'hff00, 24'hff00, 24'hff00, 24'hff00, 24'h882840, 24'hc03838, 24'hc03838, 24'hc03838, 24'he8e8f8, 24'he8e8f8, 24'hc03838, 24'hc03838, 24'hc03838, 24'h882840, 24'hff00, 24'hff00, 24'hff00, 24'h503018, 24'h885028, 24'hb8b0d0, 24'hc03838, 24'hb8b0d0, 24'hc03838, 24'hc03838, 24'hb8b0d0, 24'hc03838, 24'hb8b0d0, 24'h503018, 24'h503018, 24'hff00, 24'hff00, 24'h784040, 24'h000, 24'h882840, 24'hb8b0d0, 24'he8e8f8, 24'he8e8f8, 24'he8e8f8, 24'he8e8f8, 24'hb8b0d0, 24'h882840, 24'hd8a078, 24'h784040, 24'h000, 24'hff00, 24'hff00, 24'h503018, 24'h885028, 24'h384040, 24'h000, 24'h000, 24'h000, 24'h000, 24'h503018, 24'h885028, 24'h000, 24'h000, 24'hf8d0b8, 24'h000, 24'hff00, 24'h000, 24'hd8a078, 24'hb8b0d0, 24'h000, 24'h784040, 24'h784040, 24'h000, 24'hd8a078, 24'hd8a078, 24'hff00, 24'h000, 24'hd8a078, 24'h000, 24'hff00, 24'h000, 24'h784040, 24'hd8a078, 24'hf8d0b8, 24'hf8d0b8, 24'hf8d0b8, 24'hf8d0b8, 24'h784040, 24'h000, 24'hff00, 24'hff00, 24'h000, 24'hff00, 24'hff00, 24'h000, 24'h486060, 24'h384040, 24'h784040, 24'hd8a078, 24'hd8a078, 24'h784040, 24'h000, 24'h000, 24'hff00, 24'hff00, 24'hff00, 24'hff00, 24'hff00, 24'h000, 24'h384040, 24'h000, 24'h000, 24'h784040, 24'h784040, 24'hb8b0d0, 24'h384040, 24'h000, 24'hff00, 24'hff00, 24'hff00, 24'hff00, 24'hff00, 24'hff00, 24'h000, 24'hf8d0b8, 24'h000, 24'h000, 24'hb8b0d0, 24'h384040, 24'h384040, 24'h406888, 24'hff00, 24'hff00, 24'hff00, 24'hff00, 24'hff00, 24'hff00, 24'h000, 24'hd8a078, 24'h000, 24'h882840, 24'h384040, 24'h384040, 24'h406888, 24'h406888, 24'hff00, 24'hff00, 24'hff00, 24'hff00, 24'hff00, 24'hff00, 24'hff00, 24'hff00, 24'hff00, 24'hff00, 24'hff00, 24'h000, 24'h406888, 24'h000, 24'hff00, 24'hff00, 24'hff00, 24'hff00, 24'hff2626, 24'hff00, 24'hff00, 24'hff00, 24'hff00, 24'hff00, 24'hff00, 24'h000, 24'hc03838, 24'h000, 24'hff00, 24'hff00, 24'hff00, 24'hff2626, 24'hff9191, 24'hff2626, 24'hff00, 24'hff00, 24'hff00, 24'hff00, 24'hff00, 24'hff00, 24'h000, 24'hff00, 24'hff00, 24'hff00, 24'hff2626, 24'hff9191};
always_comb
begin
		case (keycode)
				8'h001A : 
					temp<=player_walkup[addr];// W
					 
				8'h0004 :
					temp<=player_walkleft[addr]; //A

				8'h0016 : 
					 temp<=player_walkdown[addr];// S

				8'h0007 :
					temp<=player_walkright[addr];// D
				
				default : 
					temp<=player_sit[addr];// do nothing

		endcase
end
		assign data = temp;
endmodule
