module rng(
			input [7:0] draw_x,
			input [7:0] draw_y,
			output [10:0] number
);

number = (;
endmodule
